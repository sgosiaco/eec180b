module test(
    input [3:0] SW,
    output [7:0] HEX0
);

   
   // Unit Under Test Instantiation
   seg7 UUT (SW, HEX0);



endmodule