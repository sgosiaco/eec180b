module rom_0r (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0000;
	mem[4] = 4'b0000;
	mem[5] = 4'b0000;
	mem[6] = 4'b0000;
	mem[7] = 4'b0000;
	mem[8] = 4'b0000;
	mem[9] = 4'b0000;
	mem[10] = 4'b0000;
	mem[11] = 4'b0000;
	mem[12] = 4'b0000;
	mem[13] = 4'b0000;
	mem[14] = 4'b0000;
	mem[15] = 4'b0000;
	mem[16] = 4'b0000;
	mem[17] = 4'b0000;
	mem[18] = 4'b0000;
	mem[19] = 4'b0000;
	mem[20] = 4'b0000;
	mem[21] = 4'b0000;
	mem[22] = 4'b0000;
	mem[23] = 4'b0000;
	mem[24] = 4'b0000;
	mem[25] = 4'b0000;
	mem[26] = 4'b0000;
	mem[27] = 4'b0000;
	mem[28] = 4'b0000;
	mem[29] = 4'b0000;
	mem[30] = 4'b0000;
	mem[31] = 4'b0000;
	mem[32] = 4'b0000;
	mem[33] = 4'b0000;
	mem[34] = 4'b0000;
	mem[35] = 4'b0000;
	mem[36] = 4'b0000;
	mem[37] = 4'b0000;
	mem[38] = 4'b0000;
	mem[39] = 4'b0000;
	mem[40] = 4'b0000;
	mem[41] = 4'b0000;
	mem[42] = 4'b0000;
	mem[43] = 4'b0000;
	mem[44] = 4'b0000;
	mem[45] = 4'b0000;
	mem[46] = 4'b0000;
	mem[47] = 4'b0000;
	mem[48] = 4'b0000;
	mem[49] = 4'b0000;
	mem[50] = 4'b0000;
	mem[51] = 4'b0000;
	mem[52] = 4'b0000;
	mem[53] = 4'b0000;
	mem[54] = 4'b0000;
	mem[55] = 4'b0000;
	mem[56] = 4'b0000;
	mem[57] = 4'b0000;
	mem[58] = 4'b0000;
	mem[59] = 4'b0000;
	mem[60] = 4'b0000;
	mem[61] = 4'b0000;
	mem[62] = 4'b0000;
	mem[63] = 4'b0000;
	mem[64] = 4'b0000;
	mem[65] = 4'b0000;
	mem[66] = 4'b0000;
	mem[67] = 4'b0000;
	mem[68] = 4'b0000;
	mem[69] = 4'b0000;
	mem[70] = 4'b0000;
	mem[71] = 4'b0000;
	mem[72] = 4'b0000;
	mem[73] = 4'b0000;
	mem[74] = 4'b0000;
	mem[75] = 4'b0000;
	mem[76] = 4'b0000;
	mem[77] = 4'b0000;
	mem[78] = 4'b0000;
	mem[79] = 4'b0000;
	mem[80] = 4'b0000;
	mem[81] = 4'b0000;
	mem[82] = 4'b0000;
	mem[83] = 4'b0000;
	mem[84] = 4'b0000;
	mem[85] = 4'b0000;
	mem[86] = 4'b0000;
	mem[87] = 4'b0000;
	mem[88] = 4'b0000;
	mem[89] = 4'b0000;
	mem[90] = 4'b0000;
	mem[91] = 4'b0000;
	mem[92] = 4'b0000;
	mem[93] = 4'b0000;
	mem[94] = 4'b0000;
	mem[95] = 4'b0000;
	mem[96] = 4'b0000;
	mem[97] = 4'b0000;
	mem[98] = 4'b0000;
	mem[99] = 4'b0000;
	mem[100] = 4'b0000;
	mem[101] = 4'b0000;
	mem[102] = 4'b0000;
	mem[103] = 4'b0000;
	mem[104] = 4'b0000;
	mem[105] = 4'b0000;
	mem[106] = 4'b0000;
	mem[107] = 4'b0000;
	mem[108] = 4'b0000;
	mem[109] = 4'b0000;
	mem[110] = 4'b0000;
	mem[111] = 4'b0000;
	mem[112] = 4'b0000;
	mem[113] = 4'b0000;
	mem[114] = 4'b0000;
	mem[115] = 4'b0000;
	mem[116] = 4'b0000;
	mem[117] = 4'b0000;
	mem[118] = 4'b0000;
	mem[119] = 4'b0000;
	mem[120] = 4'b0000;
	mem[121] = 4'b0000;
	mem[122] = 4'b0000;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b0000;
	mem[132] = 4'b0000;
	mem[133] = 4'b0000;
	mem[134] = 4'b0000;
	mem[135] = 4'b0000;
	mem[136] = 4'b0000;
	mem[137] = 4'b0000;
	mem[138] = 4'b0000;
	mem[139] = 4'b0000;
	mem[140] = 4'b0000;
	mem[141] = 4'b0000;
	mem[142] = 4'b0000;
	mem[143] = 4'b0000;
	mem[144] = 4'b0000;
	mem[145] = 4'b0000;
	mem[146] = 4'b0000;
	mem[147] = 4'b0000;
	mem[148] = 4'b0000;
	mem[149] = 4'b0000;
	mem[150] = 4'b0000;
	mem[151] = 4'b0000;
	mem[152] = 4'b0000;
	mem[153] = 4'b0000;
	mem[154] = 4'b0000;
	mem[155] = 4'b0000;
	mem[156] = 4'b0000;
	mem[157] = 4'b0000;
	mem[158] = 4'b0000;
	mem[159] = 4'b0000;
	mem[160] = 4'b0000;
	mem[161] = 4'b0000;
	mem[162] = 4'b0000;
	mem[163] = 4'b0000;
	mem[164] = 4'b0000;
	mem[165] = 4'b0000;
	mem[166] = 4'b0000;
	mem[167] = 4'b0000;
	mem[168] = 4'b0000;
	mem[169] = 4'b0000;
	mem[170] = 4'b0000;
	mem[171] = 4'b0000;
	mem[172] = 4'b0000;
	mem[173] = 4'b0000;
	mem[174] = 4'b0000;
	mem[175] = 4'b0000;
	mem[176] = 4'b0000;
	mem[177] = 4'b0000;
	mem[178] = 4'b0000;
	mem[179] = 4'b0000;
	mem[180] = 4'b0000;
	mem[181] = 4'b0000;
	mem[182] = 4'b0000;
	mem[183] = 4'b0000;
	mem[184] = 4'b0000;
	mem[185] = 4'b0000;
	mem[186] = 4'b0000;
	mem[187] = 4'b0000;
	mem[188] = 4'b0000;
	mem[189] = 4'b0000;
	mem[190] = 4'b0000;
	mem[191] = 4'b0000;
	mem[192] = 4'b0000;
	mem[193] = 4'b0000;
	mem[194] = 4'b0000;
	mem[195] = 4'b0000;
	mem[196] = 4'b0000;
	mem[197] = 4'b0000;
	mem[198] = 4'b0000;
	mem[199] = 4'b0000;
	mem[200] = 4'b0000;
	mem[201] = 4'b0000;
	mem[202] = 4'b0000;
	mem[203] = 4'b0000;
	mem[204] = 4'b0000;
	mem[205] = 4'b0000;
	mem[206] = 4'b0000;
	mem[207] = 4'b0000;
	mem[208] = 4'b0000;
	mem[209] = 4'b0000;
	mem[210] = 4'b0000;
	mem[211] = 4'b0000;
	mem[212] = 4'b0000;
	mem[213] = 4'b0000;
	mem[214] = 4'b0000;
	mem[215] = 4'b0000;
	mem[216] = 4'b0000;
	mem[217] = 4'b0000;
	mem[218] = 4'b0000;
	mem[219] = 4'b0000;
	mem[220] = 4'b0000;
	mem[221] = 4'b0000;
	mem[222] = 4'b0000;
	mem[223] = 4'b0000;
	mem[224] = 4'b0000;
	mem[225] = 4'b0000;
	mem[226] = 4'b0000;
	mem[227] = 4'b0000;
	mem[228] = 4'b0000;
	mem[229] = 4'b0000;
	mem[230] = 4'b0000;
	mem[231] = 4'b0000;
	mem[232] = 4'b0000;
	mem[233] = 4'b0000;
	mem[234] = 4'b0000;
	mem[235] = 4'b0000;
	mem[236] = 4'b0000;
	mem[237] = 4'b0000;
	mem[238] = 4'b0000;
	mem[239] = 4'b0000;
	mem[240] = 4'b0000;
	mem[241] = 4'b0000;
	mem[242] = 4'b0000;
	mem[243] = 4'b0000;
	mem[244] = 4'b0000;
	mem[245] = 4'b0000;
	mem[246] = 4'b0000;
	mem[247] = 4'b0000;
	mem[248] = 4'b0000;
	mem[249] = 4'b0000;
	mem[250] = 4'b0000;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0000;
	mem[260] = 4'b0000;
	mem[261] = 4'b0000;
	mem[262] = 4'b0000;
	mem[263] = 4'b0000;
	mem[264] = 4'b0000;
	mem[265] = 4'b0000;
	mem[266] = 4'b0000;
	mem[267] = 4'b0000;
	mem[268] = 4'b0000;
	mem[269] = 4'b0000;
	mem[270] = 4'b0000;
	mem[271] = 4'b0000;
	mem[272] = 4'b0000;
	mem[273] = 4'b0000;
	mem[274] = 4'b0000;
	mem[275] = 4'b0000;
	mem[276] = 4'b0000;
	mem[277] = 4'b0000;
	mem[278] = 4'b0000;
	mem[279] = 4'b0000;
	mem[280] = 4'b0000;
	mem[281] = 4'b0000;
	mem[282] = 4'b0000;
	mem[283] = 4'b0000;
	mem[284] = 4'b0000;
	mem[285] = 4'b0000;
	mem[286] = 4'b0000;
	mem[287] = 4'b0000;
	mem[288] = 4'b0000;
	mem[289] = 4'b0000;
	mem[290] = 4'b0000;
	mem[291] = 4'b0000;
	mem[292] = 4'b0000;
	mem[293] = 4'b0000;
	mem[294] = 4'b0000;
	mem[295] = 4'b0000;
	mem[296] = 4'b0000;
	mem[297] = 4'b0000;
	mem[298] = 4'b0000;
	mem[299] = 4'b0000;
	mem[300] = 4'b0000;
	mem[301] = 4'b0000;
	mem[302] = 4'b0000;
	mem[303] = 4'b0000;
	mem[304] = 4'b0000;
	mem[305] = 4'b0000;
	mem[306] = 4'b0000;
	mem[307] = 4'b0000;
	mem[308] = 4'b0000;
	mem[309] = 4'b0000;
	mem[310] = 4'b0000;
	mem[311] = 4'b0000;
	mem[312] = 4'b0000;
	mem[313] = 4'b0000;
	mem[314] = 4'b0000;
	mem[315] = 4'b0000;
	mem[316] = 4'b0000;
	mem[317] = 4'b0000;
	mem[318] = 4'b0000;
	mem[319] = 4'b0000;
	mem[320] = 4'b0000;
	mem[321] = 4'b0000;
	mem[322] = 4'b0000;
	mem[323] = 4'b0000;
	mem[324] = 4'b0000;
	mem[325] = 4'b0000;
	mem[326] = 4'b0000;
	mem[327] = 4'b0000;
	mem[328] = 4'b0000;
	mem[329] = 4'b0000;
	mem[330] = 4'b0000;
	mem[331] = 4'b0000;
	mem[332] = 4'b0000;
	mem[333] = 4'b0000;
	mem[334] = 4'b0000;
	mem[335] = 4'b0000;
	mem[336] = 4'b0000;
	mem[337] = 4'b0000;
	mem[338] = 4'b0000;
	mem[339] = 4'b0000;
	mem[340] = 4'b0000;
	mem[341] = 4'b0000;
	mem[342] = 4'b0000;
	mem[343] = 4'b0000;
	mem[344] = 4'b0000;
	mem[345] = 4'b0000;
	mem[346] = 4'b0000;
	mem[347] = 4'b0000;
	mem[348] = 4'b0000;
	mem[349] = 4'b0000;
	mem[350] = 4'b0000;
	mem[351] = 4'b0000;
	mem[352] = 4'b0000;
	mem[353] = 4'b0000;
	mem[354] = 4'b0000;
	mem[355] = 4'b0000;
	mem[356] = 4'b0000;
	mem[357] = 4'b0000;
	mem[358] = 4'b0000;
	mem[359] = 4'b0000;
	mem[360] = 4'b0000;
	mem[361] = 4'b0000;
	mem[362] = 4'b0000;
	mem[363] = 4'b0000;
	mem[364] = 4'b0000;
	mem[365] = 4'b0000;
	mem[366] = 4'b0000;
	mem[367] = 4'b0000;
	mem[368] = 4'b0000;
	mem[369] = 4'b0000;
	mem[370] = 4'b0000;
	mem[371] = 4'b0000;
	mem[372] = 4'b0000;
	mem[373] = 4'b0000;
	mem[374] = 4'b0000;
	mem[375] = 4'b0000;
	mem[376] = 4'b0000;
	mem[377] = 4'b0000;
	mem[378] = 4'b0000;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0000;
	mem[388] = 4'b0000;
	mem[389] = 4'b0000;
	mem[390] = 4'b0000;
	mem[391] = 4'b0000;
	mem[392] = 4'b0000;
	mem[393] = 4'b0000;
	mem[394] = 4'b0000;
	mem[395] = 4'b0000;
	mem[396] = 4'b0000;
	mem[397] = 4'b0000;
	mem[398] = 4'b0000;
	mem[399] = 4'b0000;
	mem[400] = 4'b0000;
	mem[401] = 4'b0000;
	mem[402] = 4'b0000;
	mem[403] = 4'b0000;
	mem[404] = 4'b0000;
	mem[405] = 4'b0000;
	mem[406] = 4'b0000;
	mem[407] = 4'b0000;
	mem[408] = 4'b0000;
	mem[409] = 4'b0000;
	mem[410] = 4'b0000;
	mem[411] = 4'b0000;
	mem[412] = 4'b0000;
	mem[413] = 4'b0000;
	mem[414] = 4'b0000;
	mem[415] = 4'b0000;
	mem[416] = 4'b0000;
	mem[417] = 4'b0000;
	mem[418] = 4'b0000;
	mem[419] = 4'b0000;
	mem[420] = 4'b0000;
	mem[421] = 4'b0000;
	mem[422] = 4'b0000;
	mem[423] = 4'b0000;
	mem[424] = 4'b0000;
	mem[425] = 4'b0000;
	mem[426] = 4'b0000;
	mem[427] = 4'b0000;
	mem[428] = 4'b0000;
	mem[429] = 4'b0000;
	mem[430] = 4'b0000;
	mem[431] = 4'b0000;
	mem[432] = 4'b0000;
	mem[433] = 4'b0000;
	mem[434] = 4'b0000;
	mem[435] = 4'b0000;
	mem[436] = 4'b0000;
	mem[437] = 4'b0000;
	mem[438] = 4'b0000;
	mem[439] = 4'b0000;
	mem[440] = 4'b0000;
	mem[441] = 4'b0000;
	mem[442] = 4'b0000;
	mem[443] = 4'b0000;
	mem[444] = 4'b0000;
	mem[445] = 4'b0000;
	mem[446] = 4'b0000;
	mem[447] = 4'b0000;
	mem[448] = 4'b0000;
	mem[449] = 4'b0000;
	mem[450] = 4'b0000;
	mem[451] = 4'b0000;
	mem[452] = 4'b0000;
	mem[453] = 4'b0000;
	mem[454] = 4'b0000;
	mem[455] = 4'b0000;
	mem[456] = 4'b0000;
	mem[457] = 4'b0000;
	mem[458] = 4'b0000;
	mem[459] = 4'b0000;
	mem[460] = 4'b0000;
	mem[461] = 4'b0000;
	mem[462] = 4'b0000;
	mem[463] = 4'b0000;
	mem[464] = 4'b0000;
	mem[465] = 4'b0000;
	mem[466] = 4'b0000;
	mem[467] = 4'b0000;
	mem[468] = 4'b0000;
	mem[469] = 4'b0000;
	mem[470] = 4'b0000;
	mem[471] = 4'b0000;
	mem[472] = 4'b0000;
	mem[473] = 4'b0000;
	mem[474] = 4'b0000;
	mem[475] = 4'b0000;
	mem[476] = 4'b0000;
	mem[477] = 4'b0000;
	mem[478] = 4'b0000;
	mem[479] = 4'b0000;
	mem[480] = 4'b0000;
	mem[481] = 4'b0000;
	mem[482] = 4'b0000;
	mem[483] = 4'b0000;
	mem[484] = 4'b0000;
	mem[485] = 4'b0000;
	mem[486] = 4'b0000;
	mem[487] = 4'b0000;
	mem[488] = 4'b0000;
	mem[489] = 4'b0000;
	mem[490] = 4'b0000;
	mem[491] = 4'b0000;
	mem[492] = 4'b0000;
	mem[493] = 4'b0000;
	mem[494] = 4'b0000;
	mem[495] = 4'b0000;
	mem[496] = 4'b0000;
	mem[497] = 4'b0000;
	mem[498] = 4'b0000;
	mem[499] = 4'b0000;
	mem[500] = 4'b0000;
	mem[501] = 4'b0000;
	mem[502] = 4'b0000;
	mem[503] = 4'b0000;
	mem[504] = 4'b0000;
	mem[505] = 4'b0000;
	mem[506] = 4'b0000;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0000;
	mem[516] = 4'b0000;
	mem[517] = 4'b0000;
	mem[518] = 4'b0000;
	mem[519] = 4'b0000;
	mem[520] = 4'b0000;
	mem[521] = 4'b0000;
	mem[522] = 4'b0000;
	mem[523] = 4'b0000;
	mem[524] = 4'b0000;
	mem[525] = 4'b0000;
	mem[526] = 4'b0000;
	mem[527] = 4'b0000;
	mem[528] = 4'b0000;
	mem[529] = 4'b0000;
	mem[530] = 4'b0000;
	mem[531] = 4'b0000;
	mem[532] = 4'b0000;
	mem[533] = 4'b0000;
	mem[534] = 4'b0000;
	mem[535] = 4'b0000;
	mem[536] = 4'b0000;
	mem[537] = 4'b0000;
	mem[538] = 4'b0000;
	mem[539] = 4'b0000;
	mem[540] = 4'b0000;
	mem[541] = 4'b0000;
	mem[542] = 4'b0000;
	mem[543] = 4'b0000;
	mem[544] = 4'b0000;
	mem[545] = 4'b0000;
	mem[546] = 4'b0000;
	mem[547] = 4'b0000;
	mem[548] = 4'b0000;
	mem[549] = 4'b0000;
	mem[550] = 4'b0000;
	mem[551] = 4'b0000;
	mem[552] = 4'b0000;
	mem[553] = 4'b0000;
	mem[554] = 4'b0000;
	mem[555] = 4'b0000;
	mem[556] = 4'b0000;
	mem[557] = 4'b0000;
	mem[558] = 4'b0000;
	mem[559] = 4'b0000;
	mem[560] = 4'b0000;
	mem[561] = 4'b0000;
	mem[562] = 4'b0000;
	mem[563] = 4'b0000;
	mem[564] = 4'b0000;
	mem[565] = 4'b0000;
	mem[566] = 4'b0000;
	mem[567] = 4'b0000;
	mem[568] = 4'b0000;
	mem[569] = 4'b0000;
	mem[570] = 4'b0000;
	mem[571] = 4'b0000;
	mem[572] = 4'b0000;
	mem[573] = 4'b0000;
	mem[574] = 4'b0000;
	mem[575] = 4'b0000;
	mem[576] = 4'b0000;
	mem[577] = 4'b0000;
	mem[578] = 4'b0000;
	mem[579] = 4'b0000;
	mem[580] = 4'b0000;
	mem[581] = 4'b0000;
	mem[582] = 4'b0000;
	mem[583] = 4'b0000;
	mem[584] = 4'b0000;
	mem[585] = 4'b0000;
	mem[586] = 4'b0000;
	mem[587] = 4'b0000;
	mem[588] = 4'b0000;
	mem[589] = 4'b0000;
	mem[590] = 4'b0000;
	mem[591] = 4'b0000;
	mem[592] = 4'b0000;
	mem[593] = 4'b0000;
	mem[594] = 4'b0000;
	mem[595] = 4'b0000;
	mem[596] = 4'b0000;
	mem[597] = 4'b0000;
	mem[598] = 4'b0000;
	mem[599] = 4'b0000;
	mem[600] = 4'b0000;
	mem[601] = 4'b0000;
	mem[602] = 4'b0000;
	mem[603] = 4'b0000;
	mem[604] = 4'b0000;
	mem[605] = 4'b0000;
	mem[606] = 4'b0000;
	mem[607] = 4'b0000;
	mem[608] = 4'b0000;
	mem[609] = 4'b0000;
	mem[610] = 4'b0000;
	mem[611] = 4'b0000;
	mem[612] = 4'b0000;
	mem[613] = 4'b0000;
	mem[614] = 4'b0000;
	mem[615] = 4'b0000;
	mem[616] = 4'b0000;
	mem[617] = 4'b0000;
	mem[618] = 4'b0000;
	mem[619] = 4'b0000;
	mem[620] = 4'b0000;
	mem[621] = 4'b0000;
	mem[622] = 4'b0000;
	mem[623] = 4'b0000;
	mem[624] = 4'b0000;
	mem[625] = 4'b0000;
	mem[626] = 4'b0000;
	mem[627] = 4'b0000;
	mem[628] = 4'b0000;
	mem[629] = 4'b0000;
	mem[630] = 4'b0000;
	mem[631] = 4'b0000;
	mem[632] = 4'b0000;
	mem[633] = 4'b0000;
	mem[634] = 4'b0000;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0000;
	mem[644] = 4'b0000;
	mem[645] = 4'b0000;
	mem[646] = 4'b0000;
	mem[647] = 4'b0000;
	mem[648] = 4'b0000;
	mem[649] = 4'b0000;
	mem[650] = 4'b0000;
	mem[651] = 4'b0000;
	mem[652] = 4'b0000;
	mem[653] = 4'b0000;
	mem[654] = 4'b0000;
	mem[655] = 4'b0000;
	mem[656] = 4'b0000;
	mem[657] = 4'b0000;
	mem[658] = 4'b0000;
	mem[659] = 4'b0000;
	mem[660] = 4'b0000;
	mem[661] = 4'b0000;
	mem[662] = 4'b0000;
	mem[663] = 4'b0000;
	mem[664] = 4'b0000;
	mem[665] = 4'b0000;
	mem[666] = 4'b0000;
	mem[667] = 4'b0000;
	mem[668] = 4'b0000;
	mem[669] = 4'b0000;
	mem[670] = 4'b0000;
	mem[671] = 4'b0000;
	mem[672] = 4'b0000;
	mem[673] = 4'b0000;
	mem[674] = 4'b0000;
	mem[675] = 4'b0000;
	mem[676] = 4'b0000;
	mem[677] = 4'b0000;
	mem[678] = 4'b0000;
	mem[679] = 4'b0000;
	mem[680] = 4'b0000;
	mem[681] = 4'b0000;
	mem[682] = 4'b0000;
	mem[683] = 4'b0000;
	mem[684] = 4'b0000;
	mem[685] = 4'b0000;
	mem[686] = 4'b0000;
	mem[687] = 4'b0000;
	mem[688] = 4'b0000;
	mem[689] = 4'b0000;
	mem[690] = 4'b0000;
	mem[691] = 4'b0000;
	mem[692] = 4'b0000;
	mem[693] = 4'b0000;
	mem[694] = 4'b0000;
	mem[695] = 4'b0000;
	mem[696] = 4'b0000;
	mem[697] = 4'b0000;
	mem[698] = 4'b0000;
	mem[699] = 4'b0000;
	mem[700] = 4'b0000;
	mem[701] = 4'b0000;
	mem[702] = 4'b0000;
	mem[703] = 4'b0000;
	mem[704] = 4'b0000;
	mem[705] = 4'b0000;
	mem[706] = 4'b0000;
	mem[707] = 4'b0000;
	mem[708] = 4'b0000;
	mem[709] = 4'b0000;
	mem[710] = 4'b0000;
	mem[711] = 4'b0000;
	mem[712] = 4'b0000;
	mem[713] = 4'b0000;
	mem[714] = 4'b0000;
	mem[715] = 4'b0000;
	mem[716] = 4'b0000;
	mem[717] = 4'b0000;
	mem[718] = 4'b0000;
	mem[719] = 4'b0000;
	mem[720] = 4'b0000;
	mem[721] = 4'b0000;
	mem[722] = 4'b0000;
	mem[723] = 4'b0000;
	mem[724] = 4'b0000;
	mem[725] = 4'b0000;
	mem[726] = 4'b0000;
	mem[727] = 4'b0000;
	mem[728] = 4'b0000;
	mem[729] = 4'b0000;
	mem[730] = 4'b0000;
	mem[731] = 4'b0000;
	mem[732] = 4'b0000;
	mem[733] = 4'b0000;
	mem[734] = 4'b0000;
	mem[735] = 4'b0000;
	mem[736] = 4'b0000;
	mem[737] = 4'b0000;
	mem[738] = 4'b0000;
	mem[739] = 4'b0000;
	mem[740] = 4'b0000;
	mem[741] = 4'b0000;
	mem[742] = 4'b0000;
	mem[743] = 4'b0000;
	mem[744] = 4'b0000;
	mem[745] = 4'b0000;
	mem[746] = 4'b0000;
	mem[747] = 4'b0000;
	mem[748] = 4'b0000;
	mem[749] = 4'b0000;
	mem[750] = 4'b0000;
	mem[751] = 4'b0000;
	mem[752] = 4'b0000;
	mem[753] = 4'b0000;
	mem[754] = 4'b0000;
	mem[755] = 4'b0000;
	mem[756] = 4'b0000;
	mem[757] = 4'b0000;
	mem[758] = 4'b0000;
	mem[759] = 4'b0000;
	mem[760] = 4'b0000;
	mem[761] = 4'b0000;
	mem[762] = 4'b0000;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0000;
	mem[772] = 4'b0000;
	mem[773] = 4'b0000;
	mem[774] = 4'b0000;
	mem[775] = 4'b0000;
	mem[776] = 4'b0000;
	mem[777] = 4'b0000;
	mem[778] = 4'b0000;
	mem[779] = 4'b0000;
	mem[780] = 4'b0000;
	mem[781] = 4'b0000;
	mem[782] = 4'b0000;
	mem[783] = 4'b0000;
	mem[784] = 4'b0000;
	mem[785] = 4'b0000;
	mem[786] = 4'b0000;
	mem[787] = 4'b0000;
	mem[788] = 4'b0000;
	mem[789] = 4'b0000;
	mem[790] = 4'b0000;
	mem[791] = 4'b0000;
	mem[792] = 4'b0000;
	mem[793] = 4'b0000;
	mem[794] = 4'b0000;
	mem[795] = 4'b0000;
	mem[796] = 4'b0000;
	mem[797] = 4'b0000;
	mem[798] = 4'b0000;
	mem[799] = 4'b0000;
	mem[800] = 4'b0000;
	mem[801] = 4'b0000;
	mem[802] = 4'b0000;
	mem[803] = 4'b0000;
	mem[804] = 4'b0000;
	mem[805] = 4'b0000;
	mem[806] = 4'b0000;
	mem[807] = 4'b0000;
	mem[808] = 4'b0000;
	mem[809] = 4'b0000;
	mem[810] = 4'b0000;
	mem[811] = 4'b0000;
	mem[812] = 4'b0000;
	mem[813] = 4'b0000;
	mem[814] = 4'b0000;
	mem[815] = 4'b0000;
	mem[816] = 4'b0000;
	mem[817] = 4'b0000;
	mem[818] = 4'b0000;
	mem[819] = 4'b0000;
	mem[820] = 4'b0000;
	mem[821] = 4'b0000;
	mem[822] = 4'b0000;
	mem[823] = 4'b0000;
	mem[824] = 4'b0000;
	mem[825] = 4'b0000;
	mem[826] = 4'b0000;
	mem[827] = 4'b0000;
	mem[828] = 4'b0000;
	mem[829] = 4'b0000;
	mem[830] = 4'b0000;
	mem[831] = 4'b0000;
	mem[832] = 4'b0000;
	mem[833] = 4'b0000;
	mem[834] = 4'b0000;
	mem[835] = 4'b0000;
	mem[836] = 4'b0000;
	mem[837] = 4'b0000;
	mem[838] = 4'b0000;
	mem[839] = 4'b0000;
	mem[840] = 4'b0000;
	mem[841] = 4'b0000;
	mem[842] = 4'b0000;
	mem[843] = 4'b0000;
	mem[844] = 4'b0000;
	mem[845] = 4'b0000;
	mem[846] = 4'b0000;
	mem[847] = 4'b0000;
	mem[848] = 4'b0000;
	mem[849] = 4'b0000;
	mem[850] = 4'b0000;
	mem[851] = 4'b0000;
	mem[852] = 4'b0000;
	mem[853] = 4'b0000;
	mem[854] = 4'b0000;
	mem[855] = 4'b0000;
	mem[856] = 4'b0000;
	mem[857] = 4'b0000;
	mem[858] = 4'b0000;
	mem[859] = 4'b0000;
	mem[860] = 4'b0000;
	mem[861] = 4'b0000;
	mem[862] = 4'b0000;
	mem[863] = 4'b0000;
	mem[864] = 4'b0000;
	mem[865] = 4'b0000;
	mem[866] = 4'b0000;
	mem[867] = 4'b0000;
	mem[868] = 4'b0000;
	mem[869] = 4'b0000;
	mem[870] = 4'b0000;
	mem[871] = 4'b0000;
	mem[872] = 4'b0000;
	mem[873] = 4'b0000;
	mem[874] = 4'b0000;
	mem[875] = 4'b0000;
	mem[876] = 4'b0000;
	mem[877] = 4'b0000;
	mem[878] = 4'b0000;
	mem[879] = 4'b0000;
	mem[880] = 4'b0000;
	mem[881] = 4'b0000;
	mem[882] = 4'b0000;
	mem[883] = 4'b0000;
	mem[884] = 4'b0000;
	mem[885] = 4'b0000;
	mem[886] = 4'b0000;
	mem[887] = 4'b0000;
	mem[888] = 4'b0000;
	mem[889] = 4'b0000;
	mem[890] = 4'b0000;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0000;
	mem[900] = 4'b0000;
	mem[901] = 4'b0000;
	mem[902] = 4'b0000;
	mem[903] = 4'b0000;
	mem[904] = 4'b0000;
	mem[905] = 4'b0000;
	mem[906] = 4'b0000;
	mem[907] = 4'b0000;
	mem[908] = 4'b0000;
	mem[909] = 4'b0000;
	mem[910] = 4'b0000;
	mem[911] = 4'b0000;
	mem[912] = 4'b0000;
	mem[913] = 4'b0000;
	mem[914] = 4'b0000;
	mem[915] = 4'b0000;
	mem[916] = 4'b0000;
	mem[917] = 4'b0000;
	mem[918] = 4'b0000;
	mem[919] = 4'b0000;
	mem[920] = 4'b0000;
	mem[921] = 4'b0000;
	mem[922] = 4'b0000;
	mem[923] = 4'b0000;
	mem[924] = 4'b0000;
	mem[925] = 4'b0000;
	mem[926] = 4'b0000;
	mem[927] = 4'b0000;
	mem[928] = 4'b0000;
	mem[929] = 4'b0000;
	mem[930] = 4'b0000;
	mem[931] = 4'b0000;
	mem[932] = 4'b0000;
	mem[933] = 4'b0000;
	mem[934] = 4'b0000;
	mem[935] = 4'b0000;
	mem[936] = 4'b0000;
	mem[937] = 4'b0000;
	mem[938] = 4'b0000;
	mem[939] = 4'b0000;
	mem[940] = 4'b0000;
	mem[941] = 4'b0000;
	mem[942] = 4'b0000;
	mem[943] = 4'b0000;
	mem[944] = 4'b0000;
	mem[945] = 4'b0000;
	mem[946] = 4'b0000;
	mem[947] = 4'b0000;
	mem[948] = 4'b0000;
	mem[949] = 4'b0000;
	mem[950] = 4'b0000;
	mem[951] = 4'b0000;
	mem[952] = 4'b0000;
	mem[953] = 4'b0000;
	mem[954] = 4'b0000;
	mem[955] = 4'b0000;
	mem[956] = 4'b0000;
	mem[957] = 4'b0000;
	mem[958] = 4'b0000;
	mem[959] = 4'b0000;
	mem[960] = 4'b0000;
	mem[961] = 4'b0000;
	mem[962] = 4'b0000;
	mem[963] = 4'b0000;
	mem[964] = 4'b0000;
	mem[965] = 4'b0000;
	mem[966] = 4'b0000;
	mem[967] = 4'b0000;
	mem[968] = 4'b0000;
	mem[969] = 4'b0000;
	mem[970] = 4'b0000;
	mem[971] = 4'b0000;
	mem[972] = 4'b0000;
	mem[973] = 4'b0000;
	mem[974] = 4'b0000;
	mem[975] = 4'b0000;
	mem[976] = 4'b0000;
	mem[977] = 4'b0000;
	mem[978] = 4'b0000;
	mem[979] = 4'b0000;
	mem[980] = 4'b0000;
	mem[981] = 4'b0000;
	mem[982] = 4'b0000;
	mem[983] = 4'b0000;
	mem[984] = 4'b0000;
	mem[985] = 4'b0000;
	mem[986] = 4'b0000;
	mem[987] = 4'b0000;
	mem[988] = 4'b0000;
	mem[989] = 4'b0000;
	mem[990] = 4'b0000;
	mem[991] = 4'b0000;
	mem[992] = 4'b0000;
	mem[993] = 4'b0000;
	mem[994] = 4'b0000;
	mem[995] = 4'b0000;
	mem[996] = 4'b0000;
	mem[997] = 4'b0000;
	mem[998] = 4'b0000;
	mem[999] = 4'b0000;
	mem[1000] = 4'b0000;
	mem[1001] = 4'b0000;
	mem[1002] = 4'b0000;
	mem[1003] = 4'b0000;
	mem[1004] = 4'b0000;
	mem[1005] = 4'b0000;
	mem[1006] = 4'b0000;
	mem[1007] = 4'b0000;
	mem[1008] = 4'b0000;
	mem[1009] = 4'b0000;
	mem[1010] = 4'b0000;
	mem[1011] = 4'b0000;
	mem[1012] = 4'b0000;
	mem[1013] = 4'b0000;
	mem[1014] = 4'b0000;
	mem[1015] = 4'b0000;
	mem[1016] = 4'b0000;
	mem[1017] = 4'b0000;
	mem[1018] = 4'b0000;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0000;
	mem[1028] = 4'b0000;
	mem[1029] = 4'b0000;
	mem[1030] = 4'b0000;
	mem[1031] = 4'b0000;
	mem[1032] = 4'b0000;
	mem[1033] = 4'b0000;
	mem[1034] = 4'b0000;
	mem[1035] = 4'b0000;
	mem[1036] = 4'b0000;
	mem[1037] = 4'b0000;
	mem[1038] = 4'b0000;
	mem[1039] = 4'b0000;
	mem[1040] = 4'b0000;
	mem[1041] = 4'b0000;
	mem[1042] = 4'b0000;
	mem[1043] = 4'b0000;
	mem[1044] = 4'b0000;
	mem[1045] = 4'b0000;
	mem[1046] = 4'b0000;
	mem[1047] = 4'b0000;
	mem[1048] = 4'b0000;
	mem[1049] = 4'b0000;
	mem[1050] = 4'b0000;
	mem[1051] = 4'b0000;
	mem[1052] = 4'b0000;
	mem[1053] = 4'b0000;
	mem[1054] = 4'b0000;
	mem[1055] = 4'b0000;
	mem[1056] = 4'b0000;
	mem[1057] = 4'b0000;
	mem[1058] = 4'b0000;
	mem[1059] = 4'b0000;
	mem[1060] = 4'b0000;
	mem[1061] = 4'b0000;
	mem[1062] = 4'b0000;
	mem[1063] = 4'b0000;
	mem[1064] = 4'b0000;
	mem[1065] = 4'b0000;
	mem[1066] = 4'b0000;
	mem[1067] = 4'b0000;
	mem[1068] = 4'b0000;
	mem[1069] = 4'b0000;
	mem[1070] = 4'b0000;
	mem[1071] = 4'b0000;
	mem[1072] = 4'b0000;
	mem[1073] = 4'b0000;
	mem[1074] = 4'b0000;
	mem[1075] = 4'b0000;
	mem[1076] = 4'b0000;
	mem[1077] = 4'b0000;
	mem[1078] = 4'b0000;
	mem[1079] = 4'b0000;
	mem[1080] = 4'b0000;
	mem[1081] = 4'b0000;
	mem[1082] = 4'b0000;
	mem[1083] = 4'b0000;
	mem[1084] = 4'b0000;
	mem[1085] = 4'b0000;
	mem[1086] = 4'b0000;
	mem[1087] = 4'b0000;
	mem[1088] = 4'b0000;
	mem[1089] = 4'b0001;
	mem[1090] = 4'b0001;
	mem[1091] = 4'b0000;
	mem[1092] = 4'b0000;
	mem[1093] = 4'b0000;
	mem[1094] = 4'b0000;
	mem[1095] = 4'b0000;
	mem[1096] = 4'b0000;
	mem[1097] = 4'b0000;
	mem[1098] = 4'b0000;
	mem[1099] = 4'b0000;
	mem[1100] = 4'b0000;
	mem[1101] = 4'b0000;
	mem[1102] = 4'b0000;
	mem[1103] = 4'b0000;
	mem[1104] = 4'b0000;
	mem[1105] = 4'b0000;
	mem[1106] = 4'b0000;
	mem[1107] = 4'b0000;
	mem[1108] = 4'b0000;
	mem[1109] = 4'b0000;
	mem[1110] = 4'b0000;
	mem[1111] = 4'b0000;
	mem[1112] = 4'b0000;
	mem[1113] = 4'b0000;
	mem[1114] = 4'b0000;
	mem[1115] = 4'b0000;
	mem[1116] = 4'b0000;
	mem[1117] = 4'b0000;
	mem[1118] = 4'b0000;
	mem[1119] = 4'b0000;
	mem[1120] = 4'b0000;
	mem[1121] = 4'b0000;
	mem[1122] = 4'b0000;
	mem[1123] = 4'b0000;
	mem[1124] = 4'b0000;
	mem[1125] = 4'b0000;
	mem[1126] = 4'b0000;
	mem[1127] = 4'b0000;
	mem[1128] = 4'b0000;
	mem[1129] = 4'b0000;
	mem[1130] = 4'b0000;
	mem[1131] = 4'b0000;
	mem[1132] = 4'b0000;
	mem[1133] = 4'b0000;
	mem[1134] = 4'b0000;
	mem[1135] = 4'b0000;
	mem[1136] = 4'b0000;
	mem[1137] = 4'b0000;
	mem[1138] = 4'b0000;
	mem[1139] = 4'b0000;
	mem[1140] = 4'b0000;
	mem[1141] = 4'b0000;
	mem[1142] = 4'b0000;
	mem[1143] = 4'b0000;
	mem[1144] = 4'b0000;
	mem[1145] = 4'b0000;
	mem[1146] = 4'b0000;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0000;
	mem[1156] = 4'b0000;
	mem[1157] = 4'b0000;
	mem[1158] = 4'b0000;
	mem[1159] = 4'b0000;
	mem[1160] = 4'b0000;
	mem[1161] = 4'b0000;
	mem[1162] = 4'b0000;
	mem[1163] = 4'b0000;
	mem[1164] = 4'b0000;
	mem[1165] = 4'b0000;
	mem[1166] = 4'b0000;
	mem[1167] = 4'b0000;
	mem[1168] = 4'b0000;
	mem[1169] = 4'b0000;
	mem[1170] = 4'b0000;
	mem[1171] = 4'b0000;
	mem[1172] = 4'b0000;
	mem[1173] = 4'b0000;
	mem[1174] = 4'b0000;
	mem[1175] = 4'b0000;
	mem[1176] = 4'b0000;
	mem[1177] = 4'b0000;
	mem[1178] = 4'b0000;
	mem[1179] = 4'b0000;
	mem[1180] = 4'b0000;
	mem[1181] = 4'b0000;
	mem[1182] = 4'b0000;
	mem[1183] = 4'b0000;
	mem[1184] = 4'b0000;
	mem[1185] = 4'b0000;
	mem[1186] = 4'b0000;
	mem[1187] = 4'b0000;
	mem[1188] = 4'b0000;
	mem[1189] = 4'b0000;
	mem[1190] = 4'b0000;
	mem[1191] = 4'b0000;
	mem[1192] = 4'b0000;
	mem[1193] = 4'b0000;
	mem[1194] = 4'b0000;
	mem[1195] = 4'b0000;
	mem[1196] = 4'b0000;
	mem[1197] = 4'b0000;
	mem[1198] = 4'b0000;
	mem[1199] = 4'b0000;
	mem[1200] = 4'b0000;
	mem[1201] = 4'b0000;
	mem[1202] = 4'b0000;
	mem[1203] = 4'b0000;
	mem[1204] = 4'b0000;
	mem[1205] = 4'b0000;
	mem[1206] = 4'b0000;
	mem[1207] = 4'b0000;
	mem[1208] = 4'b0000;
	mem[1209] = 4'b0000;
	mem[1210] = 4'b0000;
	mem[1211] = 4'b0000;
	mem[1212] = 4'b0000;
	mem[1213] = 4'b0000;
	mem[1214] = 4'b0000;
	mem[1215] = 4'b0000;
	mem[1216] = 4'b0001;
	mem[1217] = 4'b0001;
	mem[1218] = 4'b0000;
	mem[1219] = 4'b0000;
	mem[1220] = 4'b0000;
	mem[1221] = 4'b0000;
	mem[1222] = 4'b0000;
	mem[1223] = 4'b0000;
	mem[1224] = 4'b0000;
	mem[1225] = 4'b0000;
	mem[1226] = 4'b0000;
	mem[1227] = 4'b0000;
	mem[1228] = 4'b0000;
	mem[1229] = 4'b0000;
	mem[1230] = 4'b0000;
	mem[1231] = 4'b0000;
	mem[1232] = 4'b0000;
	mem[1233] = 4'b0000;
	mem[1234] = 4'b0000;
	mem[1235] = 4'b0000;
	mem[1236] = 4'b0000;
	mem[1237] = 4'b0000;
	mem[1238] = 4'b0000;
	mem[1239] = 4'b0000;
	mem[1240] = 4'b0000;
	mem[1241] = 4'b0000;
	mem[1242] = 4'b0000;
	mem[1243] = 4'b0000;
	mem[1244] = 4'b0000;
	mem[1245] = 4'b0000;
	mem[1246] = 4'b0000;
	mem[1247] = 4'b0000;
	mem[1248] = 4'b0000;
	mem[1249] = 4'b0000;
	mem[1250] = 4'b0000;
	mem[1251] = 4'b0000;
	mem[1252] = 4'b0000;
	mem[1253] = 4'b0000;
	mem[1254] = 4'b0000;
	mem[1255] = 4'b0000;
	mem[1256] = 4'b0000;
	mem[1257] = 4'b0000;
	mem[1258] = 4'b0000;
	mem[1259] = 4'b0000;
	mem[1260] = 4'b0000;
	mem[1261] = 4'b0000;
	mem[1262] = 4'b0000;
	mem[1263] = 4'b0000;
	mem[1264] = 4'b0000;
	mem[1265] = 4'b0000;
	mem[1266] = 4'b0000;
	mem[1267] = 4'b0000;
	mem[1268] = 4'b0000;
	mem[1269] = 4'b0000;
	mem[1270] = 4'b0000;
	mem[1271] = 4'b0000;
	mem[1272] = 4'b0000;
	mem[1273] = 4'b0000;
	mem[1274] = 4'b0000;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0000;
	mem[1284] = 4'b0000;
	mem[1285] = 4'b0000;
	mem[1286] = 4'b0000;
	mem[1287] = 4'b0000;
	mem[1288] = 4'b0000;
	mem[1289] = 4'b0000;
	mem[1290] = 4'b0000;
	mem[1291] = 4'b0000;
	mem[1292] = 4'b0000;
	mem[1293] = 4'b0000;
	mem[1294] = 4'b0000;
	mem[1295] = 4'b0000;
	mem[1296] = 4'b0000;
	mem[1297] = 4'b0000;
	mem[1298] = 4'b0000;
	mem[1299] = 4'b0000;
	mem[1300] = 4'b0000;
	mem[1301] = 4'b0000;
	mem[1302] = 4'b0000;
	mem[1303] = 4'b0000;
	mem[1304] = 4'b0000;
	mem[1305] = 4'b0000;
	mem[1306] = 4'b0000;
	mem[1307] = 4'b0000;
	mem[1308] = 4'b0000;
	mem[1309] = 4'b0000;
	mem[1310] = 4'b0000;
	mem[1311] = 4'b0000;
	mem[1312] = 4'b0000;
	mem[1313] = 4'b0000;
	mem[1314] = 4'b0000;
	mem[1315] = 4'b0000;
	mem[1316] = 4'b0000;
	mem[1317] = 4'b0000;
	mem[1318] = 4'b0000;
	mem[1319] = 4'b0000;
	mem[1320] = 4'b0000;
	mem[1321] = 4'b0000;
	mem[1322] = 4'b0000;
	mem[1323] = 4'b0000;
	mem[1324] = 4'b0000;
	mem[1325] = 4'b0000;
	mem[1326] = 4'b0000;
	mem[1327] = 4'b0000;
	mem[1328] = 4'b0000;
	mem[1329] = 4'b0000;
	mem[1330] = 4'b0000;
	mem[1331] = 4'b0000;
	mem[1332] = 4'b0000;
	mem[1333] = 4'b0000;
	mem[1334] = 4'b0000;
	mem[1335] = 4'b0000;
	mem[1336] = 4'b0000;
	mem[1337] = 4'b0000;
	mem[1338] = 4'b0000;
	mem[1339] = 4'b0000;
	mem[1340] = 4'b0000;
	mem[1341] = 4'b0000;
	mem[1342] = 4'b0000;
	mem[1343] = 4'b0000;
	mem[1344] = 4'b0001;
	mem[1345] = 4'b0000;
	mem[1346] = 4'b0000;
	mem[1347] = 4'b0000;
	mem[1348] = 4'b0000;
	mem[1349] = 4'b0000;
	mem[1350] = 4'b0000;
	mem[1351] = 4'b0000;
	mem[1352] = 4'b0000;
	mem[1353] = 4'b0000;
	mem[1354] = 4'b0000;
	mem[1355] = 4'b0000;
	mem[1356] = 4'b0000;
	mem[1357] = 4'b0000;
	mem[1358] = 4'b0000;
	mem[1359] = 4'b0000;
	mem[1360] = 4'b0000;
	mem[1361] = 4'b0000;
	mem[1362] = 4'b0000;
	mem[1363] = 4'b0000;
	mem[1364] = 4'b0000;
	mem[1365] = 4'b0000;
	mem[1366] = 4'b0000;
	mem[1367] = 4'b0000;
	mem[1368] = 4'b0000;
	mem[1369] = 4'b0000;
	mem[1370] = 4'b0000;
	mem[1371] = 4'b0000;
	mem[1372] = 4'b0000;
	mem[1373] = 4'b0000;
	mem[1374] = 4'b0000;
	mem[1375] = 4'b0000;
	mem[1376] = 4'b0000;
	mem[1377] = 4'b0000;
	mem[1378] = 4'b0000;
	mem[1379] = 4'b0000;
	mem[1380] = 4'b0000;
	mem[1381] = 4'b0000;
	mem[1382] = 4'b0000;
	mem[1383] = 4'b0000;
	mem[1384] = 4'b0000;
	mem[1385] = 4'b0000;
	mem[1386] = 4'b0000;
	mem[1387] = 4'b0000;
	mem[1388] = 4'b0000;
	mem[1389] = 4'b0000;
	mem[1390] = 4'b0000;
	mem[1391] = 4'b0000;
	mem[1392] = 4'b0000;
	mem[1393] = 4'b0000;
	mem[1394] = 4'b0000;
	mem[1395] = 4'b0000;
	mem[1396] = 4'b0000;
	mem[1397] = 4'b0000;
	mem[1398] = 4'b0000;
	mem[1399] = 4'b0000;
	mem[1400] = 4'b0000;
	mem[1401] = 4'b0000;
	mem[1402] = 4'b0000;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0101;
	mem[1412] = 4'b0111;
	mem[1413] = 4'b0111;
	mem[1414] = 4'b0111;
	mem[1415] = 4'b0111;
	mem[1416] = 4'b0111;
	mem[1417] = 4'b0111;
	mem[1418] = 4'b0111;
	mem[1419] = 4'b0111;
	mem[1420] = 4'b0111;
	mem[1421] = 4'b0111;
	mem[1422] = 4'b0111;
	mem[1423] = 4'b0111;
	mem[1424] = 4'b0111;
	mem[1425] = 4'b0111;
	mem[1426] = 4'b0111;
	mem[1427] = 4'b0111;
	mem[1428] = 4'b1001;
	mem[1429] = 4'b1001;
	mem[1430] = 4'b1001;
	mem[1431] = 4'b1001;
	mem[1432] = 4'b1001;
	mem[1433] = 4'b1001;
	mem[1434] = 4'b1001;
	mem[1435] = 4'b1001;
	mem[1436] = 4'b1001;
	mem[1437] = 4'b1001;
	mem[1438] = 4'b1001;
	mem[1439] = 4'b1001;
	mem[1440] = 4'b1001;
	mem[1441] = 4'b1001;
	mem[1442] = 4'b1001;
	mem[1443] = 4'b1001;
	mem[1444] = 4'b1001;
	mem[1445] = 4'b0010;
	mem[1446] = 4'b0000;
	mem[1447] = 4'b0000;
	mem[1448] = 4'b0000;
	mem[1449] = 4'b0000;
	mem[1450] = 4'b0000;
	mem[1451] = 4'b0000;
	mem[1452] = 4'b0000;
	mem[1453] = 4'b0000;
	mem[1454] = 4'b0000;
	mem[1455] = 4'b0000;
	mem[1456] = 4'b0000;
	mem[1457] = 4'b0000;
	mem[1458] = 4'b0000;
	mem[1459] = 4'b0000;
	mem[1460] = 4'b0000;
	mem[1461] = 4'b0000;
	mem[1462] = 4'b0000;
	mem[1463] = 4'b0000;
	mem[1464] = 4'b0000;
	mem[1465] = 4'b0000;
	mem[1466] = 4'b0000;
	mem[1467] = 4'b0000;
	mem[1468] = 4'b0000;
	mem[1469] = 4'b0000;
	mem[1470] = 4'b0000;
	mem[1471] = 4'b0000;
	mem[1472] = 4'b0000;
	mem[1473] = 4'b0000;
	mem[1474] = 4'b0000;
	mem[1475] = 4'b0000;
	mem[1476] = 4'b0000;
	mem[1477] = 4'b0000;
	mem[1478] = 4'b0000;
	mem[1479] = 4'b0110;
	mem[1480] = 4'b1001;
	mem[1481] = 4'b1010;
	mem[1482] = 4'b1001;
	mem[1483] = 4'b1001;
	mem[1484] = 4'b1001;
	mem[1485] = 4'b1001;
	mem[1486] = 4'b1001;
	mem[1487] = 4'b1001;
	mem[1488] = 4'b1001;
	mem[1489] = 4'b1001;
	mem[1490] = 4'b1001;
	mem[1491] = 4'b1001;
	mem[1492] = 4'b1001;
	mem[1493] = 4'b1001;
	mem[1494] = 4'b1001;
	mem[1495] = 4'b1001;
	mem[1496] = 4'b1001;
	mem[1497] = 4'b1001;
	mem[1498] = 4'b1001;
	mem[1499] = 4'b1001;
	mem[1500] = 4'b1001;
	mem[1501] = 4'b1001;
	mem[1502] = 4'b1001;
	mem[1503] = 4'b1001;
	mem[1504] = 4'b1001;
	mem[1505] = 4'b1001;
	mem[1506] = 4'b1001;
	mem[1507] = 4'b1001;
	mem[1508] = 4'b1001;
	mem[1509] = 4'b1001;
	mem[1510] = 4'b1001;
	mem[1511] = 4'b1001;
	mem[1512] = 4'b1001;
	mem[1513] = 4'b0011;
	mem[1514] = 4'b0000;
	mem[1515] = 4'b0000;
	mem[1516] = 4'b0000;
	mem[1517] = 4'b0000;
	mem[1518] = 4'b0000;
	mem[1519] = 4'b0000;
	mem[1520] = 4'b0000;
	mem[1521] = 4'b0000;
	mem[1522] = 4'b0000;
	mem[1523] = 4'b0000;
	mem[1524] = 4'b0000;
	mem[1525] = 4'b0000;
	mem[1526] = 4'b0000;
	mem[1527] = 4'b0000;
	mem[1528] = 4'b0000;
	mem[1529] = 4'b0000;
	mem[1530] = 4'b0000;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0111;
	mem[1540] = 4'b1100;
	mem[1541] = 4'b1100;
	mem[1542] = 4'b1100;
	mem[1543] = 4'b1100;
	mem[1544] = 4'b1100;
	mem[1545] = 4'b1100;
	mem[1546] = 4'b1100;
	mem[1547] = 4'b1100;
	mem[1548] = 4'b1100;
	mem[1549] = 4'b1100;
	mem[1550] = 4'b1100;
	mem[1551] = 4'b1100;
	mem[1552] = 4'b1100;
	mem[1553] = 4'b1100;
	mem[1554] = 4'b1100;
	mem[1555] = 4'b1100;
	mem[1556] = 4'b1111;
	mem[1557] = 4'b1111;
	mem[1558] = 4'b1111;
	mem[1559] = 4'b1111;
	mem[1560] = 4'b1111;
	mem[1561] = 4'b1111;
	mem[1562] = 4'b1111;
	mem[1563] = 4'b1111;
	mem[1564] = 4'b1111;
	mem[1565] = 4'b1111;
	mem[1566] = 4'b1111;
	mem[1567] = 4'b1111;
	mem[1568] = 4'b1111;
	mem[1569] = 4'b1111;
	mem[1570] = 4'b1111;
	mem[1571] = 4'b1111;
	mem[1572] = 4'b1111;
	mem[1573] = 4'b0100;
	mem[1574] = 4'b0000;
	mem[1575] = 4'b0000;
	mem[1576] = 4'b0000;
	mem[1577] = 4'b0000;
	mem[1578] = 4'b0000;
	mem[1579] = 4'b0000;
	mem[1580] = 4'b0000;
	mem[1581] = 4'b0000;
	mem[1582] = 4'b0000;
	mem[1583] = 4'b0000;
	mem[1584] = 4'b0000;
	mem[1585] = 4'b0000;
	mem[1586] = 4'b0000;
	mem[1587] = 4'b0000;
	mem[1588] = 4'b0000;
	mem[1589] = 4'b0000;
	mem[1590] = 4'b0000;
	mem[1591] = 4'b0000;
	mem[1592] = 4'b0000;
	mem[1593] = 4'b0000;
	mem[1594] = 4'b0000;
	mem[1595] = 4'b0000;
	mem[1596] = 4'b0000;
	mem[1597] = 4'b0000;
	mem[1598] = 4'b0000;
	mem[1599] = 4'b0000;
	mem[1600] = 4'b0000;
	mem[1601] = 4'b0000;
	mem[1602] = 4'b0000;
	mem[1603] = 4'b0000;
	mem[1604] = 4'b0000;
	mem[1605] = 4'b0000;
	mem[1606] = 4'b0001;
	mem[1607] = 4'b1100;
	mem[1608] = 4'b1111;
	mem[1609] = 4'b1111;
	mem[1610] = 4'b1111;
	mem[1611] = 4'b1111;
	mem[1612] = 4'b1111;
	mem[1613] = 4'b1111;
	mem[1614] = 4'b1111;
	mem[1615] = 4'b1111;
	mem[1616] = 4'b1111;
	mem[1617] = 4'b1111;
	mem[1618] = 4'b1111;
	mem[1619] = 4'b1111;
	mem[1620] = 4'b1111;
	mem[1621] = 4'b1111;
	mem[1622] = 4'b1111;
	mem[1623] = 4'b1111;
	mem[1624] = 4'b1111;
	mem[1625] = 4'b1111;
	mem[1626] = 4'b1111;
	mem[1627] = 4'b1111;
	mem[1628] = 4'b1111;
	mem[1629] = 4'b1111;
	mem[1630] = 4'b1111;
	mem[1631] = 4'b1111;
	mem[1632] = 4'b1111;
	mem[1633] = 4'b1111;
	mem[1634] = 4'b1111;
	mem[1635] = 4'b1111;
	mem[1636] = 4'b1111;
	mem[1637] = 4'b1111;
	mem[1638] = 4'b1111;
	mem[1639] = 4'b1111;
	mem[1640] = 4'b1111;
	mem[1641] = 4'b0110;
	mem[1642] = 4'b0000;
	mem[1643] = 4'b0000;
	mem[1644] = 4'b0000;
	mem[1645] = 4'b0000;
	mem[1646] = 4'b0000;
	mem[1647] = 4'b0000;
	mem[1648] = 4'b0000;
	mem[1649] = 4'b0000;
	mem[1650] = 4'b0000;
	mem[1651] = 4'b0000;
	mem[1652] = 4'b0000;
	mem[1653] = 4'b0000;
	mem[1654] = 4'b0000;
	mem[1655] = 4'b0000;
	mem[1656] = 4'b0000;
	mem[1657] = 4'b0000;
	mem[1658] = 4'b0000;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0111;
	mem[1668] = 4'b1100;
	mem[1669] = 4'b1101;
	mem[1670] = 4'b1101;
	mem[1671] = 4'b1101;
	mem[1672] = 4'b1101;
	mem[1673] = 4'b1101;
	mem[1674] = 4'b1101;
	mem[1675] = 4'b1101;
	mem[1676] = 4'b1101;
	mem[1677] = 4'b1101;
	mem[1678] = 4'b1101;
	mem[1679] = 4'b1101;
	mem[1680] = 4'b1101;
	mem[1681] = 4'b1101;
	mem[1682] = 4'b1101;
	mem[1683] = 4'b1101;
	mem[1684] = 4'b1111;
	mem[1685] = 4'b1111;
	mem[1686] = 4'b1111;
	mem[1687] = 4'b1111;
	mem[1688] = 4'b1111;
	mem[1689] = 4'b1111;
	mem[1690] = 4'b1111;
	mem[1691] = 4'b1111;
	mem[1692] = 4'b1111;
	mem[1693] = 4'b1111;
	mem[1694] = 4'b1111;
	mem[1695] = 4'b1111;
	mem[1696] = 4'b1111;
	mem[1697] = 4'b1111;
	mem[1698] = 4'b1111;
	mem[1699] = 4'b1111;
	mem[1700] = 4'b1111;
	mem[1701] = 4'b0111;
	mem[1702] = 4'b0100;
	mem[1703] = 4'b0100;
	mem[1704] = 4'b0100;
	mem[1705] = 4'b0100;
	mem[1706] = 4'b0100;
	mem[1707] = 4'b0100;
	mem[1708] = 4'b0100;
	mem[1709] = 4'b0100;
	mem[1710] = 4'b0100;
	mem[1711] = 4'b0100;
	mem[1712] = 4'b0100;
	mem[1713] = 4'b0100;
	mem[1714] = 4'b0100;
	mem[1715] = 4'b0100;
	mem[1716] = 4'b0100;
	mem[1717] = 4'b0100;
	mem[1718] = 4'b0100;
	mem[1719] = 4'b0100;
	mem[1720] = 4'b0100;
	mem[1721] = 4'b0100;
	mem[1722] = 4'b0100;
	mem[1723] = 4'b0100;
	mem[1724] = 4'b0101;
	mem[1725] = 4'b0101;
	mem[1726] = 4'b0101;
	mem[1727] = 4'b0101;
	mem[1728] = 4'b0100;
	mem[1729] = 4'b0100;
	mem[1730] = 4'b0100;
	mem[1731] = 4'b0101;
	mem[1732] = 4'b0100;
	mem[1733] = 4'b0100;
	mem[1734] = 4'b0101;
	mem[1735] = 4'b1101;
	mem[1736] = 4'b1111;
	mem[1737] = 4'b1111;
	mem[1738] = 4'b1111;
	mem[1739] = 4'b1111;
	mem[1740] = 4'b1111;
	mem[1741] = 4'b1111;
	mem[1742] = 4'b1111;
	mem[1743] = 4'b1111;
	mem[1744] = 4'b1111;
	mem[1745] = 4'b1111;
	mem[1746] = 4'b1111;
	mem[1747] = 4'b1111;
	mem[1748] = 4'b1111;
	mem[1749] = 4'b1111;
	mem[1750] = 4'b1111;
	mem[1751] = 4'b1111;
	mem[1752] = 4'b1111;
	mem[1753] = 4'b1111;
	mem[1754] = 4'b1111;
	mem[1755] = 4'b1111;
	mem[1756] = 4'b1111;
	mem[1757] = 4'b1111;
	mem[1758] = 4'b1111;
	mem[1759] = 4'b1111;
	mem[1760] = 4'b1111;
	mem[1761] = 4'b1111;
	mem[1762] = 4'b1111;
	mem[1763] = 4'b1111;
	mem[1764] = 4'b1111;
	mem[1765] = 4'b1111;
	mem[1766] = 4'b1111;
	mem[1767] = 4'b1111;
	mem[1768] = 4'b1111;
	mem[1769] = 4'b1001;
	mem[1770] = 4'b0101;
	mem[1771] = 4'b0101;
	mem[1772] = 4'b0101;
	mem[1773] = 4'b0110;
	mem[1774] = 4'b0110;
	mem[1775] = 4'b0110;
	mem[1776] = 4'b0110;
	mem[1777] = 4'b0110;
	mem[1778] = 4'b0101;
	mem[1779] = 4'b0101;
	mem[1780] = 4'b0101;
	mem[1781] = 4'b0101;
	mem[1782] = 4'b0101;
	mem[1783] = 4'b0110;
	mem[1784] = 4'b0000;
	mem[1785] = 4'b0000;
	mem[1786] = 4'b0000;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0111;
	mem[1796] = 4'b1100;
	mem[1797] = 4'b1101;
	mem[1798] = 4'b1101;
	mem[1799] = 4'b1101;
	mem[1800] = 4'b1101;
	mem[1801] = 4'b1101;
	mem[1802] = 4'b1101;
	mem[1803] = 4'b1101;
	mem[1804] = 4'b1101;
	mem[1805] = 4'b1101;
	mem[1806] = 4'b1101;
	mem[1807] = 4'b1101;
	mem[1808] = 4'b1101;
	mem[1809] = 4'b1101;
	mem[1810] = 4'b1101;
	mem[1811] = 4'b1101;
	mem[1812] = 4'b1111;
	mem[1813] = 4'b1111;
	mem[1814] = 4'b1111;
	mem[1815] = 4'b1111;
	mem[1816] = 4'b1111;
	mem[1817] = 4'b1111;
	mem[1818] = 4'b1111;
	mem[1819] = 4'b1111;
	mem[1820] = 4'b1111;
	mem[1821] = 4'b1111;
	mem[1822] = 4'b1111;
	mem[1823] = 4'b1111;
	mem[1824] = 4'b1111;
	mem[1825] = 4'b1111;
	mem[1826] = 4'b1111;
	mem[1827] = 4'b1111;
	mem[1828] = 4'b1111;
	mem[1829] = 4'b0111;
	mem[1830] = 4'b0101;
	mem[1831] = 4'b0101;
	mem[1832] = 4'b0101;
	mem[1833] = 4'b0101;
	mem[1834] = 4'b0101;
	mem[1835] = 4'b0101;
	mem[1836] = 4'b0101;
	mem[1837] = 4'b0101;
	mem[1838] = 4'b0101;
	mem[1839] = 4'b0101;
	mem[1840] = 4'b0101;
	mem[1841] = 4'b0101;
	mem[1842] = 4'b0101;
	mem[1843] = 4'b0101;
	mem[1844] = 4'b0101;
	mem[1845] = 4'b0101;
	mem[1846] = 4'b0101;
	mem[1847] = 4'b0101;
	mem[1848] = 4'b0101;
	mem[1849] = 4'b0101;
	mem[1850] = 4'b0101;
	mem[1851] = 4'b0101;
	mem[1852] = 4'b0101;
	mem[1853] = 4'b0101;
	mem[1854] = 4'b0101;
	mem[1855] = 4'b0101;
	mem[1856] = 4'b0110;
	mem[1857] = 4'b0101;
	mem[1858] = 4'b0101;
	mem[1859] = 4'b0101;
	mem[1860] = 4'b0101;
	mem[1861] = 4'b0110;
	mem[1862] = 4'b0110;
	mem[1863] = 4'b1101;
	mem[1864] = 4'b1111;
	mem[1865] = 4'b1111;
	mem[1866] = 4'b1111;
	mem[1867] = 4'b1111;
	mem[1868] = 4'b1111;
	mem[1869] = 4'b1111;
	mem[1870] = 4'b1111;
	mem[1871] = 4'b1111;
	mem[1872] = 4'b1111;
	mem[1873] = 4'b1111;
	mem[1874] = 4'b1111;
	mem[1875] = 4'b1111;
	mem[1876] = 4'b1111;
	mem[1877] = 4'b1111;
	mem[1878] = 4'b1111;
	mem[1879] = 4'b1111;
	mem[1880] = 4'b1111;
	mem[1881] = 4'b1111;
	mem[1882] = 4'b1111;
	mem[1883] = 4'b1111;
	mem[1884] = 4'b1111;
	mem[1885] = 4'b1111;
	mem[1886] = 4'b1111;
	mem[1887] = 4'b1111;
	mem[1888] = 4'b1111;
	mem[1889] = 4'b1111;
	mem[1890] = 4'b1111;
	mem[1891] = 4'b1111;
	mem[1892] = 4'b1111;
	mem[1893] = 4'b1111;
	mem[1894] = 4'b1111;
	mem[1895] = 4'b1111;
	mem[1896] = 4'b1111;
	mem[1897] = 4'b1001;
	mem[1898] = 4'b0110;
	mem[1899] = 4'b0110;
	mem[1900] = 4'b0110;
	mem[1901] = 4'b0111;
	mem[1902] = 4'b0111;
	mem[1903] = 4'b0110;
	mem[1904] = 4'b0110;
	mem[1905] = 4'b0111;
	mem[1906] = 4'b0111;
	mem[1907] = 4'b0110;
	mem[1908] = 4'b0110;
	mem[1909] = 4'b0110;
	mem[1910] = 4'b0110;
	mem[1911] = 4'b0110;
	mem[1912] = 4'b0000;
	mem[1913] = 4'b0000;
	mem[1914] = 4'b0000;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0111;
	mem[1924] = 4'b1100;
	mem[1925] = 4'b1101;
	mem[1926] = 4'b1101;
	mem[1927] = 4'b1101;
	mem[1928] = 4'b1101;
	mem[1929] = 4'b1101;
	mem[1930] = 4'b1101;
	mem[1931] = 4'b1101;
	mem[1932] = 4'b1101;
	mem[1933] = 4'b1101;
	mem[1934] = 4'b1101;
	mem[1935] = 4'b1101;
	mem[1936] = 4'b1101;
	mem[1937] = 4'b1101;
	mem[1938] = 4'b1101;
	mem[1939] = 4'b1101;
	mem[1940] = 4'b1111;
	mem[1941] = 4'b1111;
	mem[1942] = 4'b1111;
	mem[1943] = 4'b1111;
	mem[1944] = 4'b1111;
	mem[1945] = 4'b1111;
	mem[1946] = 4'b1111;
	mem[1947] = 4'b1111;
	mem[1948] = 4'b1111;
	mem[1949] = 4'b1111;
	mem[1950] = 4'b1111;
	mem[1951] = 4'b1111;
	mem[1952] = 4'b1111;
	mem[1953] = 4'b1111;
	mem[1954] = 4'b1111;
	mem[1955] = 4'b1111;
	mem[1956] = 4'b1111;
	mem[1957] = 4'b0111;
	mem[1958] = 4'b0101;
	mem[1959] = 4'b0101;
	mem[1960] = 4'b0101;
	mem[1961] = 4'b0101;
	mem[1962] = 4'b0101;
	mem[1963] = 4'b0101;
	mem[1964] = 4'b0101;
	mem[1965] = 4'b0101;
	mem[1966] = 4'b0101;
	mem[1967] = 4'b0101;
	mem[1968] = 4'b0101;
	mem[1969] = 4'b0101;
	mem[1970] = 4'b0101;
	mem[1971] = 4'b0101;
	mem[1972] = 4'b0101;
	mem[1973] = 4'b0101;
	mem[1974] = 4'b0101;
	mem[1975] = 4'b0101;
	mem[1976] = 4'b0101;
	mem[1977] = 4'b0101;
	mem[1978] = 4'b0101;
	mem[1979] = 4'b0101;
	mem[1980] = 4'b0101;
	mem[1981] = 4'b0101;
	mem[1982] = 4'b0101;
	mem[1983] = 4'b0101;
	mem[1984] = 4'b0101;
	mem[1985] = 4'b0110;
	mem[1986] = 4'b0110;
	mem[1987] = 4'b0110;
	mem[1988] = 4'b0110;
	mem[1989] = 4'b0110;
	mem[1990] = 4'b0110;
	mem[1991] = 4'b1101;
	mem[1992] = 4'b1111;
	mem[1993] = 4'b1111;
	mem[1994] = 4'b1111;
	mem[1995] = 4'b1111;
	mem[1996] = 4'b1111;
	mem[1997] = 4'b1111;
	mem[1998] = 4'b1111;
	mem[1999] = 4'b1111;
	mem[2000] = 4'b1111;
	mem[2001] = 4'b1111;
	mem[2002] = 4'b1111;
	mem[2003] = 4'b1111;
	mem[2004] = 4'b1111;
	mem[2005] = 4'b1111;
	mem[2006] = 4'b1111;
	mem[2007] = 4'b1111;
	mem[2008] = 4'b1111;
	mem[2009] = 4'b1111;
	mem[2010] = 4'b1111;
	mem[2011] = 4'b1111;
	mem[2012] = 4'b1111;
	mem[2013] = 4'b1111;
	mem[2014] = 4'b1111;
	mem[2015] = 4'b1111;
	mem[2016] = 4'b1111;
	mem[2017] = 4'b1111;
	mem[2018] = 4'b1111;
	mem[2019] = 4'b1111;
	mem[2020] = 4'b1111;
	mem[2021] = 4'b1111;
	mem[2022] = 4'b1111;
	mem[2023] = 4'b1111;
	mem[2024] = 4'b1111;
	mem[2025] = 4'b1001;
	mem[2026] = 4'b0110;
	mem[2027] = 4'b0110;
	mem[2028] = 4'b0111;
	mem[2029] = 4'b0111;
	mem[2030] = 4'b0110;
	mem[2031] = 4'b0110;
	mem[2032] = 4'b0110;
	mem[2033] = 4'b0110;
	mem[2034] = 4'b0110;
	mem[2035] = 4'b0111;
	mem[2036] = 4'b0110;
	mem[2037] = 4'b0110;
	mem[2038] = 4'b0110;
	mem[2039] = 4'b0110;
	mem[2040] = 4'b0000;
	mem[2041] = 4'b0000;
	mem[2042] = 4'b0000;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0111;
	mem[2052] = 4'b1100;
	mem[2053] = 4'b1101;
	mem[2054] = 4'b1101;
	mem[2055] = 4'b1101;
	mem[2056] = 4'b1101;
	mem[2057] = 4'b1101;
	mem[2058] = 4'b1101;
	mem[2059] = 4'b1101;
	mem[2060] = 4'b1101;
	mem[2061] = 4'b1101;
	mem[2062] = 4'b1101;
	mem[2063] = 4'b1101;
	mem[2064] = 4'b1101;
	mem[2065] = 4'b1101;
	mem[2066] = 4'b1101;
	mem[2067] = 4'b1101;
	mem[2068] = 4'b1111;
	mem[2069] = 4'b1111;
	mem[2070] = 4'b1111;
	mem[2071] = 4'b1111;
	mem[2072] = 4'b1111;
	mem[2073] = 4'b1111;
	mem[2074] = 4'b1111;
	mem[2075] = 4'b1111;
	mem[2076] = 4'b1111;
	mem[2077] = 4'b1111;
	mem[2078] = 4'b1111;
	mem[2079] = 4'b1111;
	mem[2080] = 4'b1111;
	mem[2081] = 4'b1111;
	mem[2082] = 4'b1111;
	mem[2083] = 4'b1111;
	mem[2084] = 4'b1111;
	mem[2085] = 4'b0111;
	mem[2086] = 4'b0101;
	mem[2087] = 4'b0101;
	mem[2088] = 4'b0101;
	mem[2089] = 4'b0101;
	mem[2090] = 4'b0101;
	mem[2091] = 4'b0101;
	mem[2092] = 4'b0101;
	mem[2093] = 4'b0101;
	mem[2094] = 4'b0101;
	mem[2095] = 4'b0101;
	mem[2096] = 4'b0101;
	mem[2097] = 4'b0101;
	mem[2098] = 4'b0101;
	mem[2099] = 4'b0101;
	mem[2100] = 4'b0101;
	mem[2101] = 4'b0101;
	mem[2102] = 4'b0101;
	mem[2103] = 4'b0101;
	mem[2104] = 4'b0101;
	mem[2105] = 4'b0101;
	mem[2106] = 4'b0110;
	mem[2107] = 4'b0110;
	mem[2108] = 4'b0110;
	mem[2109] = 4'b0101;
	mem[2110] = 4'b0101;
	mem[2111] = 4'b0101;
	mem[2112] = 4'b0110;
	mem[2113] = 4'b0101;
	mem[2114] = 4'b0110;
	mem[2115] = 4'b0110;
	mem[2116] = 4'b0110;
	mem[2117] = 4'b0110;
	mem[2118] = 4'b0110;
	mem[2119] = 4'b1101;
	mem[2120] = 4'b1111;
	mem[2121] = 4'b1111;
	mem[2122] = 4'b1111;
	mem[2123] = 4'b1111;
	mem[2124] = 4'b1111;
	mem[2125] = 4'b1111;
	mem[2126] = 4'b1111;
	mem[2127] = 4'b1111;
	mem[2128] = 4'b1111;
	mem[2129] = 4'b1111;
	mem[2130] = 4'b1111;
	mem[2131] = 4'b1111;
	mem[2132] = 4'b1111;
	mem[2133] = 4'b1111;
	mem[2134] = 4'b1111;
	mem[2135] = 4'b1111;
	mem[2136] = 4'b1111;
	mem[2137] = 4'b1111;
	mem[2138] = 4'b1111;
	mem[2139] = 4'b1111;
	mem[2140] = 4'b1111;
	mem[2141] = 4'b1111;
	mem[2142] = 4'b1111;
	mem[2143] = 4'b1111;
	mem[2144] = 4'b1111;
	mem[2145] = 4'b1111;
	mem[2146] = 4'b1111;
	mem[2147] = 4'b1111;
	mem[2148] = 4'b1111;
	mem[2149] = 4'b1111;
	mem[2150] = 4'b1111;
	mem[2151] = 4'b1111;
	mem[2152] = 4'b1111;
	mem[2153] = 4'b1001;
	mem[2154] = 4'b0110;
	mem[2155] = 4'b0110;
	mem[2156] = 4'b0111;
	mem[2157] = 4'b0111;
	mem[2158] = 4'b0110;
	mem[2159] = 4'b0110;
	mem[2160] = 4'b0110;
	mem[2161] = 4'b0111;
	mem[2162] = 4'b0111;
	mem[2163] = 4'b0111;
	mem[2164] = 4'b0111;
	mem[2165] = 4'b0110;
	mem[2166] = 4'b0110;
	mem[2167] = 4'b0110;
	mem[2168] = 4'b0000;
	mem[2169] = 4'b0000;
	mem[2170] = 4'b0000;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0111;
	mem[2180] = 4'b1100;
	mem[2181] = 4'b1101;
	mem[2182] = 4'b1101;
	mem[2183] = 4'b1101;
	mem[2184] = 4'b1101;
	mem[2185] = 4'b1101;
	mem[2186] = 4'b1101;
	mem[2187] = 4'b1101;
	mem[2188] = 4'b1101;
	mem[2189] = 4'b1101;
	mem[2190] = 4'b1101;
	mem[2191] = 4'b1101;
	mem[2192] = 4'b1101;
	mem[2193] = 4'b1101;
	mem[2194] = 4'b1101;
	mem[2195] = 4'b1101;
	mem[2196] = 4'b1111;
	mem[2197] = 4'b1111;
	mem[2198] = 4'b1111;
	mem[2199] = 4'b1111;
	mem[2200] = 4'b1111;
	mem[2201] = 4'b1111;
	mem[2202] = 4'b1111;
	mem[2203] = 4'b1111;
	mem[2204] = 4'b1111;
	mem[2205] = 4'b1111;
	mem[2206] = 4'b1111;
	mem[2207] = 4'b1111;
	mem[2208] = 4'b1111;
	mem[2209] = 4'b1111;
	mem[2210] = 4'b1111;
	mem[2211] = 4'b1111;
	mem[2212] = 4'b1111;
	mem[2213] = 4'b0111;
	mem[2214] = 4'b0101;
	mem[2215] = 4'b0101;
	mem[2216] = 4'b0101;
	mem[2217] = 4'b0101;
	mem[2218] = 4'b0101;
	mem[2219] = 4'b0101;
	mem[2220] = 4'b0101;
	mem[2221] = 4'b0101;
	mem[2222] = 4'b0101;
	mem[2223] = 4'b0101;
	mem[2224] = 4'b0101;
	mem[2225] = 4'b0101;
	mem[2226] = 4'b0101;
	mem[2227] = 4'b0101;
	mem[2228] = 4'b0101;
	mem[2229] = 4'b0101;
	mem[2230] = 4'b0101;
	mem[2231] = 4'b0101;
	mem[2232] = 4'b0101;
	mem[2233] = 4'b0110;
	mem[2234] = 4'b0110;
	mem[2235] = 4'b0101;
	mem[2236] = 4'b0101;
	mem[2237] = 4'b0110;
	mem[2238] = 4'b0101;
	mem[2239] = 4'b0101;
	mem[2240] = 4'b0110;
	mem[2241] = 4'b0110;
	mem[2242] = 4'b0101;
	mem[2243] = 4'b0101;
	mem[2244] = 4'b0110;
	mem[2245] = 4'b0110;
	mem[2246] = 4'b0110;
	mem[2247] = 4'b1101;
	mem[2248] = 4'b1111;
	mem[2249] = 4'b1111;
	mem[2250] = 4'b1111;
	mem[2251] = 4'b1111;
	mem[2252] = 4'b1111;
	mem[2253] = 4'b1111;
	mem[2254] = 4'b1111;
	mem[2255] = 4'b1111;
	mem[2256] = 4'b1111;
	mem[2257] = 4'b1111;
	mem[2258] = 4'b1111;
	mem[2259] = 4'b1111;
	mem[2260] = 4'b1111;
	mem[2261] = 4'b1111;
	mem[2262] = 4'b1111;
	mem[2263] = 4'b1111;
	mem[2264] = 4'b1111;
	mem[2265] = 4'b1111;
	mem[2266] = 4'b1111;
	mem[2267] = 4'b1111;
	mem[2268] = 4'b1111;
	mem[2269] = 4'b1111;
	mem[2270] = 4'b1111;
	mem[2271] = 4'b1111;
	mem[2272] = 4'b1111;
	mem[2273] = 4'b1111;
	mem[2274] = 4'b1111;
	mem[2275] = 4'b1111;
	mem[2276] = 4'b1111;
	mem[2277] = 4'b1111;
	mem[2278] = 4'b1111;
	mem[2279] = 4'b1111;
	mem[2280] = 4'b1111;
	mem[2281] = 4'b1001;
	mem[2282] = 4'b0110;
	mem[2283] = 4'b0110;
	mem[2284] = 4'b0110;
	mem[2285] = 4'b0111;
	mem[2286] = 4'b0110;
	mem[2287] = 4'b0111;
	mem[2288] = 4'b0111;
	mem[2289] = 4'b0111;
	mem[2290] = 4'b0111;
	mem[2291] = 4'b0111;
	mem[2292] = 4'b0111;
	mem[2293] = 4'b0110;
	mem[2294] = 4'b0110;
	mem[2295] = 4'b0110;
	mem[2296] = 4'b0000;
	mem[2297] = 4'b0000;
	mem[2298] = 4'b0000;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0111;
	mem[2308] = 4'b1100;
	mem[2309] = 4'b1101;
	mem[2310] = 4'b1101;
	mem[2311] = 4'b1101;
	mem[2312] = 4'b1101;
	mem[2313] = 4'b1101;
	mem[2314] = 4'b1101;
	mem[2315] = 4'b1101;
	mem[2316] = 4'b1101;
	mem[2317] = 4'b1101;
	mem[2318] = 4'b1101;
	mem[2319] = 4'b1101;
	mem[2320] = 4'b1101;
	mem[2321] = 4'b1101;
	mem[2322] = 4'b1101;
	mem[2323] = 4'b1101;
	mem[2324] = 4'b1111;
	mem[2325] = 4'b1111;
	mem[2326] = 4'b1111;
	mem[2327] = 4'b1111;
	mem[2328] = 4'b1111;
	mem[2329] = 4'b1111;
	mem[2330] = 4'b1111;
	mem[2331] = 4'b1111;
	mem[2332] = 4'b1111;
	mem[2333] = 4'b1111;
	mem[2334] = 4'b1111;
	mem[2335] = 4'b1111;
	mem[2336] = 4'b1111;
	mem[2337] = 4'b1111;
	mem[2338] = 4'b1111;
	mem[2339] = 4'b1111;
	mem[2340] = 4'b1111;
	mem[2341] = 4'b0111;
	mem[2342] = 4'b0101;
	mem[2343] = 4'b0101;
	mem[2344] = 4'b0101;
	mem[2345] = 4'b0101;
	mem[2346] = 4'b0101;
	mem[2347] = 4'b0101;
	mem[2348] = 4'b0101;
	mem[2349] = 4'b0101;
	mem[2350] = 4'b0101;
	mem[2351] = 4'b0101;
	mem[2352] = 4'b0101;
	mem[2353] = 4'b0101;
	mem[2354] = 4'b0101;
	mem[2355] = 4'b0101;
	mem[2356] = 4'b0101;
	mem[2357] = 4'b0101;
	mem[2358] = 4'b0101;
	mem[2359] = 4'b0101;
	mem[2360] = 4'b0101;
	mem[2361] = 4'b0101;
	mem[2362] = 4'b0110;
	mem[2363] = 4'b0101;
	mem[2364] = 4'b0101;
	mem[2365] = 4'b0101;
	mem[2366] = 4'b0110;
	mem[2367] = 4'b0101;
	mem[2368] = 4'b0101;
	mem[2369] = 4'b0110;
	mem[2370] = 4'b0110;
	mem[2371] = 4'b0110;
	mem[2372] = 4'b0110;
	mem[2373] = 4'b0110;
	mem[2374] = 4'b0110;
	mem[2375] = 4'b1101;
	mem[2376] = 4'b1111;
	mem[2377] = 4'b1111;
	mem[2378] = 4'b1111;
	mem[2379] = 4'b1111;
	mem[2380] = 4'b1111;
	mem[2381] = 4'b1111;
	mem[2382] = 4'b1111;
	mem[2383] = 4'b1111;
	mem[2384] = 4'b1111;
	mem[2385] = 4'b1111;
	mem[2386] = 4'b1111;
	mem[2387] = 4'b1111;
	mem[2388] = 4'b1111;
	mem[2389] = 4'b1111;
	mem[2390] = 4'b1111;
	mem[2391] = 4'b1111;
	mem[2392] = 4'b1111;
	mem[2393] = 4'b1111;
	mem[2394] = 4'b1111;
	mem[2395] = 4'b1111;
	mem[2396] = 4'b1111;
	mem[2397] = 4'b1111;
	mem[2398] = 4'b1111;
	mem[2399] = 4'b1111;
	mem[2400] = 4'b1111;
	mem[2401] = 4'b1111;
	mem[2402] = 4'b1111;
	mem[2403] = 4'b1111;
	mem[2404] = 4'b1111;
	mem[2405] = 4'b1111;
	mem[2406] = 4'b1111;
	mem[2407] = 4'b1111;
	mem[2408] = 4'b1111;
	mem[2409] = 4'b1001;
	mem[2410] = 4'b0110;
	mem[2411] = 4'b0110;
	mem[2412] = 4'b0110;
	mem[2413] = 4'b0111;
	mem[2414] = 4'b0111;
	mem[2415] = 4'b0111;
	mem[2416] = 4'b0111;
	mem[2417] = 4'b0111;
	mem[2418] = 4'b0111;
	mem[2419] = 4'b0111;
	mem[2420] = 4'b0111;
	mem[2421] = 4'b0110;
	mem[2422] = 4'b0110;
	mem[2423] = 4'b0110;
	mem[2424] = 4'b0000;
	mem[2425] = 4'b0000;
	mem[2426] = 4'b0001;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0111;
	mem[2436] = 4'b1100;
	mem[2437] = 4'b1101;
	mem[2438] = 4'b1101;
	mem[2439] = 4'b1101;
	mem[2440] = 4'b1101;
	mem[2441] = 4'b1101;
	mem[2442] = 4'b1101;
	mem[2443] = 4'b1101;
	mem[2444] = 4'b1101;
	mem[2445] = 4'b1101;
	mem[2446] = 4'b1101;
	mem[2447] = 4'b1101;
	mem[2448] = 4'b1101;
	mem[2449] = 4'b1101;
	mem[2450] = 4'b1101;
	mem[2451] = 4'b1101;
	mem[2452] = 4'b1111;
	mem[2453] = 4'b1111;
	mem[2454] = 4'b1111;
	mem[2455] = 4'b1111;
	mem[2456] = 4'b1111;
	mem[2457] = 4'b1111;
	mem[2458] = 4'b1111;
	mem[2459] = 4'b1111;
	mem[2460] = 4'b1111;
	mem[2461] = 4'b1111;
	mem[2462] = 4'b1111;
	mem[2463] = 4'b1111;
	mem[2464] = 4'b1111;
	mem[2465] = 4'b1111;
	mem[2466] = 4'b1111;
	mem[2467] = 4'b1111;
	mem[2468] = 4'b1111;
	mem[2469] = 4'b1000;
	mem[2470] = 4'b0101;
	mem[2471] = 4'b0101;
	mem[2472] = 4'b0101;
	mem[2473] = 4'b0101;
	mem[2474] = 4'b0101;
	mem[2475] = 4'b0101;
	mem[2476] = 4'b0101;
	mem[2477] = 4'b0101;
	mem[2478] = 4'b0101;
	mem[2479] = 4'b0101;
	mem[2480] = 4'b0101;
	mem[2481] = 4'b0101;
	mem[2482] = 4'b0101;
	mem[2483] = 4'b0101;
	mem[2484] = 4'b0101;
	mem[2485] = 4'b0101;
	mem[2486] = 4'b0101;
	mem[2487] = 4'b0110;
	mem[2488] = 4'b0101;
	mem[2489] = 4'b0101;
	mem[2490] = 4'b0101;
	mem[2491] = 4'b0110;
	mem[2492] = 4'b0101;
	mem[2493] = 4'b0101;
	mem[2494] = 4'b0110;
	mem[2495] = 4'b0110;
	mem[2496] = 4'b0110;
	mem[2497] = 4'b0110;
	mem[2498] = 4'b0110;
	mem[2499] = 4'b0110;
	mem[2500] = 4'b0110;
	mem[2501] = 4'b0110;
	mem[2502] = 4'b0110;
	mem[2503] = 4'b1101;
	mem[2504] = 4'b1111;
	mem[2505] = 4'b1111;
	mem[2506] = 4'b1111;
	mem[2507] = 4'b1111;
	mem[2508] = 4'b1111;
	mem[2509] = 4'b1111;
	mem[2510] = 4'b1111;
	mem[2511] = 4'b1111;
	mem[2512] = 4'b1111;
	mem[2513] = 4'b1111;
	mem[2514] = 4'b1111;
	mem[2515] = 4'b1111;
	mem[2516] = 4'b1111;
	mem[2517] = 4'b1111;
	mem[2518] = 4'b1111;
	mem[2519] = 4'b1111;
	mem[2520] = 4'b1111;
	mem[2521] = 4'b1111;
	mem[2522] = 4'b1111;
	mem[2523] = 4'b1111;
	mem[2524] = 4'b1111;
	mem[2525] = 4'b1111;
	mem[2526] = 4'b1111;
	mem[2527] = 4'b1111;
	mem[2528] = 4'b1111;
	mem[2529] = 4'b1111;
	mem[2530] = 4'b1111;
	mem[2531] = 4'b1111;
	mem[2532] = 4'b1111;
	mem[2533] = 4'b1111;
	mem[2534] = 4'b1111;
	mem[2535] = 4'b1111;
	mem[2536] = 4'b1111;
	mem[2537] = 4'b1001;
	mem[2538] = 4'b0110;
	mem[2539] = 4'b0110;
	mem[2540] = 4'b0110;
	mem[2541] = 4'b0110;
	mem[2542] = 4'b0111;
	mem[2543] = 4'b0111;
	mem[2544] = 4'b0111;
	mem[2545] = 4'b0111;
	mem[2546] = 4'b0111;
	mem[2547] = 4'b0111;
	mem[2548] = 4'b0111;
	mem[2549] = 4'b0110;
	mem[2550] = 4'b0110;
	mem[2551] = 4'b0111;
	mem[2552] = 4'b0001;
	mem[2553] = 4'b0001;
	mem[2554] = 4'b0000;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b0111;
	mem[2564] = 4'b1100;
	mem[2565] = 4'b1101;
	mem[2566] = 4'b1101;
	mem[2567] = 4'b1101;
	mem[2568] = 4'b1101;
	mem[2569] = 4'b1101;
	mem[2570] = 4'b1101;
	mem[2571] = 4'b1101;
	mem[2572] = 4'b1101;
	mem[2573] = 4'b1101;
	mem[2574] = 4'b1101;
	mem[2575] = 4'b1101;
	mem[2576] = 4'b1101;
	mem[2577] = 4'b1101;
	mem[2578] = 4'b1101;
	mem[2579] = 4'b1101;
	mem[2580] = 4'b1111;
	mem[2581] = 4'b1111;
	mem[2582] = 4'b1111;
	mem[2583] = 4'b1111;
	mem[2584] = 4'b1111;
	mem[2585] = 4'b1111;
	mem[2586] = 4'b1111;
	mem[2587] = 4'b1111;
	mem[2588] = 4'b1111;
	mem[2589] = 4'b1111;
	mem[2590] = 4'b1111;
	mem[2591] = 4'b1111;
	mem[2592] = 4'b1111;
	mem[2593] = 4'b1111;
	mem[2594] = 4'b1111;
	mem[2595] = 4'b1111;
	mem[2596] = 4'b1111;
	mem[2597] = 4'b1000;
	mem[2598] = 4'b0101;
	mem[2599] = 4'b0101;
	mem[2600] = 4'b0101;
	mem[2601] = 4'b0101;
	mem[2602] = 4'b0101;
	mem[2603] = 4'b0101;
	mem[2604] = 4'b0101;
	mem[2605] = 4'b0101;
	mem[2606] = 4'b0101;
	mem[2607] = 4'b0101;
	mem[2608] = 4'b0101;
	mem[2609] = 4'b0101;
	mem[2610] = 4'b0101;
	mem[2611] = 4'b0101;
	mem[2612] = 4'b0101;
	mem[2613] = 4'b0101;
	mem[2614] = 4'b0101;
	mem[2615] = 4'b0101;
	mem[2616] = 4'b0110;
	mem[2617] = 4'b0101;
	mem[2618] = 4'b0101;
	mem[2619] = 4'b0110;
	mem[2620] = 4'b0110;
	mem[2621] = 4'b0101;
	mem[2622] = 4'b0110;
	mem[2623] = 4'b0110;
	mem[2624] = 4'b0110;
	mem[2625] = 4'b0110;
	mem[2626] = 4'b0110;
	mem[2627] = 4'b0110;
	mem[2628] = 4'b0110;
	mem[2629] = 4'b0110;
	mem[2630] = 4'b0110;
	mem[2631] = 4'b1101;
	mem[2632] = 4'b1111;
	mem[2633] = 4'b1111;
	mem[2634] = 4'b1111;
	mem[2635] = 4'b1111;
	mem[2636] = 4'b1111;
	mem[2637] = 4'b1111;
	mem[2638] = 4'b1111;
	mem[2639] = 4'b1111;
	mem[2640] = 4'b1111;
	mem[2641] = 4'b1111;
	mem[2642] = 4'b1111;
	mem[2643] = 4'b1111;
	mem[2644] = 4'b1111;
	mem[2645] = 4'b1111;
	mem[2646] = 4'b1111;
	mem[2647] = 4'b1111;
	mem[2648] = 4'b1111;
	mem[2649] = 4'b1111;
	mem[2650] = 4'b1111;
	mem[2651] = 4'b1111;
	mem[2652] = 4'b1111;
	mem[2653] = 4'b1111;
	mem[2654] = 4'b1111;
	mem[2655] = 4'b1111;
	mem[2656] = 4'b1111;
	mem[2657] = 4'b1111;
	mem[2658] = 4'b1111;
	mem[2659] = 4'b1111;
	mem[2660] = 4'b1111;
	mem[2661] = 4'b1111;
	mem[2662] = 4'b1111;
	mem[2663] = 4'b1111;
	mem[2664] = 4'b1111;
	mem[2665] = 4'b1010;
	mem[2666] = 4'b0110;
	mem[2667] = 4'b0110;
	mem[2668] = 4'b0110;
	mem[2669] = 4'b0110;
	mem[2670] = 4'b0110;
	mem[2671] = 4'b0111;
	mem[2672] = 4'b0111;
	mem[2673] = 4'b0111;
	mem[2674] = 4'b0111;
	mem[2675] = 4'b0111;
	mem[2676] = 4'b0110;
	mem[2677] = 4'b0110;
	mem[2678] = 4'b0110;
	mem[2679] = 4'b1000;
	mem[2680] = 4'b0000;
	mem[2681] = 4'b0000;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b0111;
	mem[2692] = 4'b1100;
	mem[2693] = 4'b1101;
	mem[2694] = 4'b1101;
	mem[2695] = 4'b1101;
	mem[2696] = 4'b1101;
	mem[2697] = 4'b1101;
	mem[2698] = 4'b1101;
	mem[2699] = 4'b1101;
	mem[2700] = 4'b1101;
	mem[2701] = 4'b1101;
	mem[2702] = 4'b1101;
	mem[2703] = 4'b1101;
	mem[2704] = 4'b1101;
	mem[2705] = 4'b1101;
	mem[2706] = 4'b1101;
	mem[2707] = 4'b1101;
	mem[2708] = 4'b1111;
	mem[2709] = 4'b1111;
	mem[2710] = 4'b1111;
	mem[2711] = 4'b1111;
	mem[2712] = 4'b1111;
	mem[2713] = 4'b1111;
	mem[2714] = 4'b1111;
	mem[2715] = 4'b1111;
	mem[2716] = 4'b1111;
	mem[2717] = 4'b1111;
	mem[2718] = 4'b1111;
	mem[2719] = 4'b1111;
	mem[2720] = 4'b1111;
	mem[2721] = 4'b1111;
	mem[2722] = 4'b1111;
	mem[2723] = 4'b1111;
	mem[2724] = 4'b1111;
	mem[2725] = 4'b1000;
	mem[2726] = 4'b0101;
	mem[2727] = 4'b0101;
	mem[2728] = 4'b0101;
	mem[2729] = 4'b0101;
	mem[2730] = 4'b0101;
	mem[2731] = 4'b0101;
	mem[2732] = 4'b0101;
	mem[2733] = 4'b0101;
	mem[2734] = 4'b0101;
	mem[2735] = 4'b0101;
	mem[2736] = 4'b0101;
	mem[2737] = 4'b0101;
	mem[2738] = 4'b0101;
	mem[2739] = 4'b0101;
	mem[2740] = 4'b0101;
	mem[2741] = 4'b0101;
	mem[2742] = 4'b0110;
	mem[2743] = 4'b0101;
	mem[2744] = 4'b0101;
	mem[2745] = 4'b0110;
	mem[2746] = 4'b0101;
	mem[2747] = 4'b0101;
	mem[2748] = 4'b0110;
	mem[2749] = 4'b0110;
	mem[2750] = 4'b0110;
	mem[2751] = 4'b0110;
	mem[2752] = 4'b0110;
	mem[2753] = 4'b0110;
	mem[2754] = 4'b0110;
	mem[2755] = 4'b0110;
	mem[2756] = 4'b0110;
	mem[2757] = 4'b0110;
	mem[2758] = 4'b0110;
	mem[2759] = 4'b1101;
	mem[2760] = 4'b1111;
	mem[2761] = 4'b1111;
	mem[2762] = 4'b1111;
	mem[2763] = 4'b1111;
	mem[2764] = 4'b1111;
	mem[2765] = 4'b1111;
	mem[2766] = 4'b1111;
	mem[2767] = 4'b1111;
	mem[2768] = 4'b1111;
	mem[2769] = 4'b1111;
	mem[2770] = 4'b1111;
	mem[2771] = 4'b1111;
	mem[2772] = 4'b1111;
	mem[2773] = 4'b1111;
	mem[2774] = 4'b1111;
	mem[2775] = 4'b1111;
	mem[2776] = 4'b1111;
	mem[2777] = 4'b1111;
	mem[2778] = 4'b1111;
	mem[2779] = 4'b1111;
	mem[2780] = 4'b1111;
	mem[2781] = 4'b1111;
	mem[2782] = 4'b1111;
	mem[2783] = 4'b1111;
	mem[2784] = 4'b1111;
	mem[2785] = 4'b1111;
	mem[2786] = 4'b1111;
	mem[2787] = 4'b1110;
	mem[2788] = 4'b1111;
	mem[2789] = 4'b1111;
	mem[2790] = 4'b1111;
	mem[2791] = 4'b1111;
	mem[2792] = 4'b1111;
	mem[2793] = 4'b1010;
	mem[2794] = 4'b0111;
	mem[2795] = 4'b0110;
	mem[2796] = 4'b0110;
	mem[2797] = 4'b0110;
	mem[2798] = 4'b0110;
	mem[2799] = 4'b0110;
	mem[2800] = 4'b0110;
	mem[2801] = 4'b0110;
	mem[2802] = 4'b0110;
	mem[2803] = 4'b0110;
	mem[2804] = 4'b0110;
	mem[2805] = 4'b0110;
	mem[2806] = 4'b0111;
	mem[2807] = 4'b1000;
	mem[2808] = 4'b0000;
	mem[2809] = 4'b0000;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b0111;
	mem[2820] = 4'b1100;
	mem[2821] = 4'b1101;
	mem[2822] = 4'b1101;
	mem[2823] = 4'b1101;
	mem[2824] = 4'b1101;
	mem[2825] = 4'b1101;
	mem[2826] = 4'b1101;
	mem[2827] = 4'b1101;
	mem[2828] = 4'b1101;
	mem[2829] = 4'b1101;
	mem[2830] = 4'b1101;
	mem[2831] = 4'b1101;
	mem[2832] = 4'b1101;
	mem[2833] = 4'b1101;
	mem[2834] = 4'b1101;
	mem[2835] = 4'b1101;
	mem[2836] = 4'b1111;
	mem[2837] = 4'b1111;
	mem[2838] = 4'b1111;
	mem[2839] = 4'b1111;
	mem[2840] = 4'b1111;
	mem[2841] = 4'b1111;
	mem[2842] = 4'b1111;
	mem[2843] = 4'b1111;
	mem[2844] = 4'b1111;
	mem[2845] = 4'b1111;
	mem[2846] = 4'b1111;
	mem[2847] = 4'b1111;
	mem[2848] = 4'b1111;
	mem[2849] = 4'b1111;
	mem[2850] = 4'b1111;
	mem[2851] = 4'b1111;
	mem[2852] = 4'b1111;
	mem[2853] = 4'b1000;
	mem[2854] = 4'b0101;
	mem[2855] = 4'b0101;
	mem[2856] = 4'b0101;
	mem[2857] = 4'b0101;
	mem[2858] = 4'b0101;
	mem[2859] = 4'b0101;
	mem[2860] = 4'b0101;
	mem[2861] = 4'b0101;
	mem[2862] = 4'b0101;
	mem[2863] = 4'b0101;
	mem[2864] = 4'b0101;
	mem[2865] = 4'b0101;
	mem[2866] = 4'b0101;
	mem[2867] = 4'b0101;
	mem[2868] = 4'b0101;
	mem[2869] = 4'b0101;
	mem[2870] = 4'b0101;
	mem[2871] = 4'b0110;
	mem[2872] = 4'b0110;
	mem[2873] = 4'b0110;
	mem[2874] = 4'b0110;
	mem[2875] = 4'b0101;
	mem[2876] = 4'b0101;
	mem[2877] = 4'b0110;
	mem[2878] = 4'b0110;
	mem[2879] = 4'b0110;
	mem[2880] = 4'b0110;
	mem[2881] = 4'b0110;
	mem[2882] = 4'b0110;
	mem[2883] = 4'b0110;
	mem[2884] = 4'b0110;
	mem[2885] = 4'b0110;
	mem[2886] = 4'b0110;
	mem[2887] = 4'b1101;
	mem[2888] = 4'b1111;
	mem[2889] = 4'b1111;
	mem[2890] = 4'b1111;
	mem[2891] = 4'b1111;
	mem[2892] = 4'b1111;
	mem[2893] = 4'b1111;
	mem[2894] = 4'b1111;
	mem[2895] = 4'b1111;
	mem[2896] = 4'b1111;
	mem[2897] = 4'b1111;
	mem[2898] = 4'b1111;
	mem[2899] = 4'b1111;
	mem[2900] = 4'b1111;
	mem[2901] = 4'b1111;
	mem[2902] = 4'b1111;
	mem[2903] = 4'b1111;
	mem[2904] = 4'b1111;
	mem[2905] = 4'b1111;
	mem[2906] = 4'b1111;
	mem[2907] = 4'b1111;
	mem[2908] = 4'b1111;
	mem[2909] = 4'b1111;
	mem[2910] = 4'b1111;
	mem[2911] = 4'b1111;
	mem[2912] = 4'b1111;
	mem[2913] = 4'b1110;
	mem[2914] = 4'b1101;
	mem[2915] = 4'b1101;
	mem[2916] = 4'b1101;
	mem[2917] = 4'b1101;
	mem[2918] = 4'b1110;
	mem[2919] = 4'b1111;
	mem[2920] = 4'b1111;
	mem[2921] = 4'b1010;
	mem[2922] = 4'b0111;
	mem[2923] = 4'b0111;
	mem[2924] = 4'b0110;
	mem[2925] = 4'b0110;
	mem[2926] = 4'b0110;
	mem[2927] = 4'b0110;
	mem[2928] = 4'b0110;
	mem[2929] = 4'b0110;
	mem[2930] = 4'b0110;
	mem[2931] = 4'b0110;
	mem[2932] = 4'b0110;
	mem[2933] = 4'b0110;
	mem[2934] = 4'b1000;
	mem[2935] = 4'b0111;
	mem[2936] = 4'b0000;
	mem[2937] = 4'b0000;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b0111;
	mem[2948] = 4'b1100;
	mem[2949] = 4'b1101;
	mem[2950] = 4'b1101;
	mem[2951] = 4'b1101;
	mem[2952] = 4'b1101;
	mem[2953] = 4'b1101;
	mem[2954] = 4'b1101;
	mem[2955] = 4'b1101;
	mem[2956] = 4'b1101;
	mem[2957] = 4'b1101;
	mem[2958] = 4'b1101;
	mem[2959] = 4'b1101;
	mem[2960] = 4'b1101;
	mem[2961] = 4'b1101;
	mem[2962] = 4'b1101;
	mem[2963] = 4'b1101;
	mem[2964] = 4'b1111;
	mem[2965] = 4'b1111;
	mem[2966] = 4'b1111;
	mem[2967] = 4'b1111;
	mem[2968] = 4'b1111;
	mem[2969] = 4'b1111;
	mem[2970] = 4'b1111;
	mem[2971] = 4'b1111;
	mem[2972] = 4'b1111;
	mem[2973] = 4'b1111;
	mem[2974] = 4'b1111;
	mem[2975] = 4'b1111;
	mem[2976] = 4'b1111;
	mem[2977] = 4'b1111;
	mem[2978] = 4'b1111;
	mem[2979] = 4'b1111;
	mem[2980] = 4'b1111;
	mem[2981] = 4'b1000;
	mem[2982] = 4'b0101;
	mem[2983] = 4'b0101;
	mem[2984] = 4'b0101;
	mem[2985] = 4'b0101;
	mem[2986] = 4'b0101;
	mem[2987] = 4'b0101;
	mem[2988] = 4'b0101;
	mem[2989] = 4'b0101;
	mem[2990] = 4'b0101;
	mem[2991] = 4'b0101;
	mem[2992] = 4'b0101;
	mem[2993] = 4'b0101;
	mem[2994] = 4'b0110;
	mem[2995] = 4'b0110;
	mem[2996] = 4'b0110;
	mem[2997] = 4'b0101;
	mem[2998] = 4'b0101;
	mem[2999] = 4'b0101;
	mem[3000] = 4'b0110;
	mem[3001] = 4'b0110;
	mem[3002] = 4'b0110;
	mem[3003] = 4'b0110;
	mem[3004] = 4'b0110;
	mem[3005] = 4'b0110;
	mem[3006] = 4'b0110;
	mem[3007] = 4'b0110;
	mem[3008] = 4'b0110;
	mem[3009] = 4'b0110;
	mem[3010] = 4'b0110;
	mem[3011] = 4'b0110;
	mem[3012] = 4'b0110;
	mem[3013] = 4'b0110;
	mem[3014] = 4'b0110;
	mem[3015] = 4'b1101;
	mem[3016] = 4'b1111;
	mem[3017] = 4'b1111;
	mem[3018] = 4'b1111;
	mem[3019] = 4'b1111;
	mem[3020] = 4'b1111;
	mem[3021] = 4'b1111;
	mem[3022] = 4'b1111;
	mem[3023] = 4'b1111;
	mem[3024] = 4'b1111;
	mem[3025] = 4'b1111;
	mem[3026] = 4'b1111;
	mem[3027] = 4'b1111;
	mem[3028] = 4'b1111;
	mem[3029] = 4'b1111;
	mem[3030] = 4'b1111;
	mem[3031] = 4'b1111;
	mem[3032] = 4'b1111;
	mem[3033] = 4'b1111;
	mem[3034] = 4'b1111;
	mem[3035] = 4'b1111;
	mem[3036] = 4'b1111;
	mem[3037] = 4'b1111;
	mem[3038] = 4'b1111;
	mem[3039] = 4'b1111;
	mem[3040] = 4'b1110;
	mem[3041] = 4'b1101;
	mem[3042] = 4'b1101;
	mem[3043] = 4'b1101;
	mem[3044] = 4'b1101;
	mem[3045] = 4'b1101;
	mem[3046] = 4'b1101;
	mem[3047] = 4'b1110;
	mem[3048] = 4'b1111;
	mem[3049] = 4'b1010;
	mem[3050] = 4'b0111;
	mem[3051] = 4'b0111;
	mem[3052] = 4'b0111;
	mem[3053] = 4'b0110;
	mem[3054] = 4'b0110;
	mem[3055] = 4'b0110;
	mem[3056] = 4'b0110;
	mem[3057] = 4'b0110;
	mem[3058] = 4'b0110;
	mem[3059] = 4'b0110;
	mem[3060] = 4'b0110;
	mem[3061] = 4'b0111;
	mem[3062] = 4'b1000;
	mem[3063] = 4'b0111;
	mem[3064] = 4'b0000;
	mem[3065] = 4'b0000;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b0111;
	mem[3076] = 4'b1100;
	mem[3077] = 4'b1101;
	mem[3078] = 4'b1101;
	mem[3079] = 4'b1101;
	mem[3080] = 4'b1101;
	mem[3081] = 4'b1101;
	mem[3082] = 4'b1101;
	mem[3083] = 4'b1101;
	mem[3084] = 4'b1101;
	mem[3085] = 4'b1101;
	mem[3086] = 4'b1101;
	mem[3087] = 4'b1101;
	mem[3088] = 4'b1101;
	mem[3089] = 4'b1101;
	mem[3090] = 4'b1101;
	mem[3091] = 4'b1101;
	mem[3092] = 4'b1111;
	mem[3093] = 4'b1111;
	mem[3094] = 4'b1111;
	mem[3095] = 4'b1111;
	mem[3096] = 4'b1111;
	mem[3097] = 4'b1111;
	mem[3098] = 4'b1111;
	mem[3099] = 4'b1111;
	mem[3100] = 4'b1111;
	mem[3101] = 4'b1111;
	mem[3102] = 4'b1111;
	mem[3103] = 4'b1111;
	mem[3104] = 4'b1111;
	mem[3105] = 4'b1111;
	mem[3106] = 4'b1111;
	mem[3107] = 4'b1111;
	mem[3108] = 4'b1111;
	mem[3109] = 4'b1000;
	mem[3110] = 4'b0101;
	mem[3111] = 4'b0101;
	mem[3112] = 4'b0101;
	mem[3113] = 4'b0101;
	mem[3114] = 4'b0101;
	mem[3115] = 4'b0101;
	mem[3116] = 4'b0101;
	mem[3117] = 4'b0101;
	mem[3118] = 4'b0101;
	mem[3119] = 4'b0101;
	mem[3120] = 4'b0101;
	mem[3121] = 4'b0101;
	mem[3122] = 4'b0110;
	mem[3123] = 4'b0110;
	mem[3124] = 4'b0101;
	mem[3125] = 4'b0101;
	mem[3126] = 4'b0110;
	mem[3127] = 4'b0101;
	mem[3128] = 4'b0101;
	mem[3129] = 4'b0110;
	mem[3130] = 4'b0110;
	mem[3131] = 4'b0110;
	mem[3132] = 4'b0110;
	mem[3133] = 4'b0110;
	mem[3134] = 4'b0110;
	mem[3135] = 4'b0110;
	mem[3136] = 4'b0110;
	mem[3137] = 4'b0110;
	mem[3138] = 4'b0110;
	mem[3139] = 4'b0110;
	mem[3140] = 4'b0110;
	mem[3141] = 4'b0110;
	mem[3142] = 4'b0110;
	mem[3143] = 4'b1101;
	mem[3144] = 4'b1111;
	mem[3145] = 4'b1111;
	mem[3146] = 4'b1111;
	mem[3147] = 4'b1111;
	mem[3148] = 4'b1111;
	mem[3149] = 4'b1111;
	mem[3150] = 4'b1111;
	mem[3151] = 4'b1111;
	mem[3152] = 4'b1111;
	mem[3153] = 4'b1111;
	mem[3154] = 4'b1111;
	mem[3155] = 4'b1111;
	mem[3156] = 4'b1111;
	mem[3157] = 4'b1111;
	mem[3158] = 4'b1111;
	mem[3159] = 4'b1111;
	mem[3160] = 4'b1111;
	mem[3161] = 4'b1111;
	mem[3162] = 4'b1111;
	mem[3163] = 4'b1111;
	mem[3164] = 4'b1111;
	mem[3165] = 4'b1111;
	mem[3166] = 4'b1111;
	mem[3167] = 4'b1110;
	mem[3168] = 4'b1101;
	mem[3169] = 4'b1101;
	mem[3170] = 4'b1101;
	mem[3171] = 4'b1101;
	mem[3172] = 4'b1101;
	mem[3173] = 4'b1101;
	mem[3174] = 4'b1101;
	mem[3175] = 4'b1101;
	mem[3176] = 4'b1110;
	mem[3177] = 4'b1010;
	mem[3178] = 4'b0111;
	mem[3179] = 4'b0111;
	mem[3180] = 4'b0111;
	mem[3181] = 4'b0111;
	mem[3182] = 4'b0111;
	mem[3183] = 4'b0110;
	mem[3184] = 4'b0110;
	mem[3185] = 4'b0110;
	mem[3186] = 4'b0110;
	mem[3187] = 4'b0111;
	mem[3188] = 4'b1000;
	mem[3189] = 4'b1000;
	mem[3190] = 4'b0111;
	mem[3191] = 4'b0111;
	mem[3192] = 4'b0000;
	mem[3193] = 4'b0000;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b0111;
	mem[3204] = 4'b1100;
	mem[3205] = 4'b1101;
	mem[3206] = 4'b1101;
	mem[3207] = 4'b1101;
	mem[3208] = 4'b1101;
	mem[3209] = 4'b1101;
	mem[3210] = 4'b1101;
	mem[3211] = 4'b1101;
	mem[3212] = 4'b1101;
	mem[3213] = 4'b1101;
	mem[3214] = 4'b1101;
	mem[3215] = 4'b1101;
	mem[3216] = 4'b1101;
	mem[3217] = 4'b1101;
	mem[3218] = 4'b1101;
	mem[3219] = 4'b1101;
	mem[3220] = 4'b1111;
	mem[3221] = 4'b1111;
	mem[3222] = 4'b1111;
	mem[3223] = 4'b1111;
	mem[3224] = 4'b1111;
	mem[3225] = 4'b1111;
	mem[3226] = 4'b1111;
	mem[3227] = 4'b1111;
	mem[3228] = 4'b1111;
	mem[3229] = 4'b1111;
	mem[3230] = 4'b1111;
	mem[3231] = 4'b1111;
	mem[3232] = 4'b1111;
	mem[3233] = 4'b1111;
	mem[3234] = 4'b1111;
	mem[3235] = 4'b1111;
	mem[3236] = 4'b1111;
	mem[3237] = 4'b1000;
	mem[3238] = 4'b0101;
	mem[3239] = 4'b0101;
	mem[3240] = 4'b0101;
	mem[3241] = 4'b0101;
	mem[3242] = 4'b0101;
	mem[3243] = 4'b0101;
	mem[3244] = 4'b0101;
	mem[3245] = 4'b0101;
	mem[3246] = 4'b0101;
	mem[3247] = 4'b0101;
	mem[3248] = 4'b0101;
	mem[3249] = 4'b0101;
	mem[3250] = 4'b0110;
	mem[3251] = 4'b0110;
	mem[3252] = 4'b0101;
	mem[3253] = 4'b0110;
	mem[3254] = 4'b0110;
	mem[3255] = 4'b0101;
	mem[3256] = 4'b0101;
	mem[3257] = 4'b0101;
	mem[3258] = 4'b0110;
	mem[3259] = 4'b0110;
	mem[3260] = 4'b0110;
	mem[3261] = 4'b0110;
	mem[3262] = 4'b0110;
	mem[3263] = 4'b0110;
	mem[3264] = 4'b0110;
	mem[3265] = 4'b0110;
	mem[3266] = 4'b0110;
	mem[3267] = 4'b0110;
	mem[3268] = 4'b0110;
	mem[3269] = 4'b0110;
	mem[3270] = 4'b0110;
	mem[3271] = 4'b1101;
	mem[3272] = 4'b1111;
	mem[3273] = 4'b1111;
	mem[3274] = 4'b1111;
	mem[3275] = 4'b1111;
	mem[3276] = 4'b1111;
	mem[3277] = 4'b1111;
	mem[3278] = 4'b1111;
	mem[3279] = 4'b1111;
	mem[3280] = 4'b1111;
	mem[3281] = 4'b1111;
	mem[3282] = 4'b1111;
	mem[3283] = 4'b1111;
	mem[3284] = 4'b1111;
	mem[3285] = 4'b1111;
	mem[3286] = 4'b1111;
	mem[3287] = 4'b1111;
	mem[3288] = 4'b1111;
	mem[3289] = 4'b1111;
	mem[3290] = 4'b1111;
	mem[3291] = 4'b1111;
	mem[3292] = 4'b1111;
	mem[3293] = 4'b1111;
	mem[3294] = 4'b1111;
	mem[3295] = 4'b1101;
	mem[3296] = 4'b1101;
	mem[3297] = 4'b1110;
	mem[3298] = 4'b1110;
	mem[3299] = 4'b1110;
	mem[3300] = 4'b1110;
	mem[3301] = 4'b1101;
	mem[3302] = 4'b1101;
	mem[3303] = 4'b1101;
	mem[3304] = 4'b1101;
	mem[3305] = 4'b1001;
	mem[3306] = 4'b0111;
	mem[3307] = 4'b0111;
	mem[3308] = 4'b0111;
	mem[3309] = 4'b0111;
	mem[3310] = 4'b0111;
	mem[3311] = 4'b0111;
	mem[3312] = 4'b0111;
	mem[3313] = 4'b1000;
	mem[3314] = 4'b1000;
	mem[3315] = 4'b1000;
	mem[3316] = 4'b0111;
	mem[3317] = 4'b0111;
	mem[3318] = 4'b0111;
	mem[3319] = 4'b0111;
	mem[3320] = 4'b0000;
	mem[3321] = 4'b0000;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b0111;
	mem[3332] = 4'b1100;
	mem[3333] = 4'b1101;
	mem[3334] = 4'b1101;
	mem[3335] = 4'b1101;
	mem[3336] = 4'b1101;
	mem[3337] = 4'b1101;
	mem[3338] = 4'b1101;
	mem[3339] = 4'b1101;
	mem[3340] = 4'b1101;
	mem[3341] = 4'b1101;
	mem[3342] = 4'b1101;
	mem[3343] = 4'b1101;
	mem[3344] = 4'b1101;
	mem[3345] = 4'b1101;
	mem[3346] = 4'b1101;
	mem[3347] = 4'b1101;
	mem[3348] = 4'b1111;
	mem[3349] = 4'b1111;
	mem[3350] = 4'b1111;
	mem[3351] = 4'b1111;
	mem[3352] = 4'b1111;
	mem[3353] = 4'b1111;
	mem[3354] = 4'b1111;
	mem[3355] = 4'b1111;
	mem[3356] = 4'b1111;
	mem[3357] = 4'b1111;
	mem[3358] = 4'b1111;
	mem[3359] = 4'b1111;
	mem[3360] = 4'b1111;
	mem[3361] = 4'b1111;
	mem[3362] = 4'b1111;
	mem[3363] = 4'b1111;
	mem[3364] = 4'b1111;
	mem[3365] = 4'b1000;
	mem[3366] = 4'b0101;
	mem[3367] = 4'b0101;
	mem[3368] = 4'b0101;
	mem[3369] = 4'b0101;
	mem[3370] = 4'b0101;
	mem[3371] = 4'b0101;
	mem[3372] = 4'b0101;
	mem[3373] = 4'b0101;
	mem[3374] = 4'b0101;
	mem[3375] = 4'b0101;
	mem[3376] = 4'b0110;
	mem[3377] = 4'b0110;
	mem[3378] = 4'b0110;
	mem[3379] = 4'b0101;
	mem[3380] = 4'b0110;
	mem[3381] = 4'b0110;
	mem[3382] = 4'b0110;
	mem[3383] = 4'b0101;
	mem[3384] = 4'b0101;
	mem[3385] = 4'b0110;
	mem[3386] = 4'b0111;
	mem[3387] = 4'b0110;
	mem[3388] = 4'b0110;
	mem[3389] = 4'b0110;
	mem[3390] = 4'b0110;
	mem[3391] = 4'b0110;
	mem[3392] = 4'b0110;
	mem[3393] = 4'b0110;
	mem[3394] = 4'b0110;
	mem[3395] = 4'b0110;
	mem[3396] = 4'b0110;
	mem[3397] = 4'b0110;
	mem[3398] = 4'b0110;
	mem[3399] = 4'b1101;
	mem[3400] = 4'b1111;
	mem[3401] = 4'b1111;
	mem[3402] = 4'b1111;
	mem[3403] = 4'b1111;
	mem[3404] = 4'b1111;
	mem[3405] = 4'b1111;
	mem[3406] = 4'b1111;
	mem[3407] = 4'b1111;
	mem[3408] = 4'b1111;
	mem[3409] = 4'b1111;
	mem[3410] = 4'b1111;
	mem[3411] = 4'b1111;
	mem[3412] = 4'b1111;
	mem[3413] = 4'b1111;
	mem[3414] = 4'b1111;
	mem[3415] = 4'b1111;
	mem[3416] = 4'b1111;
	mem[3417] = 4'b1111;
	mem[3418] = 4'b1111;
	mem[3419] = 4'b1111;
	mem[3420] = 4'b1111;
	mem[3421] = 4'b1111;
	mem[3422] = 4'b1111;
	mem[3423] = 4'b1101;
	mem[3424] = 4'b1101;
	mem[3425] = 4'b1111;
	mem[3426] = 4'b1111;
	mem[3427] = 4'b1111;
	mem[3428] = 4'b1111;
	mem[3429] = 4'b1110;
	mem[3430] = 4'b1101;
	mem[3431] = 4'b1101;
	mem[3432] = 4'b1101;
	mem[3433] = 4'b1001;
	mem[3434] = 4'b0111;
	mem[3435] = 4'b0111;
	mem[3436] = 4'b0111;
	mem[3437] = 4'b0111;
	mem[3438] = 4'b0111;
	mem[3439] = 4'b0111;
	mem[3440] = 4'b0111;
	mem[3441] = 4'b0111;
	mem[3442] = 4'b0111;
	mem[3443] = 4'b0111;
	mem[3444] = 4'b0111;
	mem[3445] = 4'b0111;
	mem[3446] = 4'b0111;
	mem[3447] = 4'b0111;
	mem[3448] = 4'b0000;
	mem[3449] = 4'b0000;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b0111;
	mem[3460] = 4'b1100;
	mem[3461] = 4'b1101;
	mem[3462] = 4'b1101;
	mem[3463] = 4'b1101;
	mem[3464] = 4'b1101;
	mem[3465] = 4'b1101;
	mem[3466] = 4'b1101;
	mem[3467] = 4'b1101;
	mem[3468] = 4'b1101;
	mem[3469] = 4'b1101;
	mem[3470] = 4'b1101;
	mem[3471] = 4'b1101;
	mem[3472] = 4'b1101;
	mem[3473] = 4'b1101;
	mem[3474] = 4'b1101;
	mem[3475] = 4'b1101;
	mem[3476] = 4'b1111;
	mem[3477] = 4'b1111;
	mem[3478] = 4'b1111;
	mem[3479] = 4'b1111;
	mem[3480] = 4'b1111;
	mem[3481] = 4'b1111;
	mem[3482] = 4'b1111;
	mem[3483] = 4'b1111;
	mem[3484] = 4'b1111;
	mem[3485] = 4'b1111;
	mem[3486] = 4'b1111;
	mem[3487] = 4'b1111;
	mem[3488] = 4'b1111;
	mem[3489] = 4'b1111;
	mem[3490] = 4'b1111;
	mem[3491] = 4'b1111;
	mem[3492] = 4'b1111;
	mem[3493] = 4'b1000;
	mem[3494] = 4'b0101;
	mem[3495] = 4'b0101;
	mem[3496] = 4'b0101;
	mem[3497] = 4'b0101;
	mem[3498] = 4'b0101;
	mem[3499] = 4'b0101;
	mem[3500] = 4'b0101;
	mem[3501] = 4'b0101;
	mem[3502] = 4'b0101;
	mem[3503] = 4'b0101;
	mem[3504] = 4'b0101;
	mem[3505] = 4'b0110;
	mem[3506] = 4'b0110;
	mem[3507] = 4'b0101;
	mem[3508] = 4'b0101;
	mem[3509] = 4'b0110;
	mem[3510] = 4'b0101;
	mem[3511] = 4'b0101;
	mem[3512] = 4'b0110;
	mem[3513] = 4'b0110;
	mem[3514] = 4'b0110;
	mem[3515] = 4'b0110;
	mem[3516] = 4'b0110;
	mem[3517] = 4'b0110;
	mem[3518] = 4'b0110;
	mem[3519] = 4'b0110;
	mem[3520] = 4'b0110;
	mem[3521] = 4'b0110;
	mem[3522] = 4'b0110;
	mem[3523] = 4'b0110;
	mem[3524] = 4'b0110;
	mem[3525] = 4'b0110;
	mem[3526] = 4'b0110;
	mem[3527] = 4'b1101;
	mem[3528] = 4'b1111;
	mem[3529] = 4'b1111;
	mem[3530] = 4'b1111;
	mem[3531] = 4'b1111;
	mem[3532] = 4'b1111;
	mem[3533] = 4'b1111;
	mem[3534] = 4'b1111;
	mem[3535] = 4'b1111;
	mem[3536] = 4'b1111;
	mem[3537] = 4'b1111;
	mem[3538] = 4'b1111;
	mem[3539] = 4'b1111;
	mem[3540] = 4'b1111;
	mem[3541] = 4'b1111;
	mem[3542] = 4'b1111;
	mem[3543] = 4'b1111;
	mem[3544] = 4'b1111;
	mem[3545] = 4'b1111;
	mem[3546] = 4'b1111;
	mem[3547] = 4'b1111;
	mem[3548] = 4'b1110;
	mem[3549] = 4'b1110;
	mem[3550] = 4'b1110;
	mem[3551] = 4'b1101;
	mem[3552] = 4'b1110;
	mem[3553] = 4'b1111;
	mem[3554] = 4'b1111;
	mem[3555] = 4'b1111;
	mem[3556] = 4'b1111;
	mem[3557] = 4'b1111;
	mem[3558] = 4'b1110;
	mem[3559] = 4'b1101;
	mem[3560] = 4'b1101;
	mem[3561] = 4'b1001;
	mem[3562] = 4'b0110;
	mem[3563] = 4'b0111;
	mem[3564] = 4'b0111;
	mem[3565] = 4'b0111;
	mem[3566] = 4'b0111;
	mem[3567] = 4'b0111;
	mem[3568] = 4'b0111;
	mem[3569] = 4'b0111;
	mem[3570] = 4'b0111;
	mem[3571] = 4'b0111;
	mem[3572] = 4'b0111;
	mem[3573] = 4'b0111;
	mem[3574] = 4'b0111;
	mem[3575] = 4'b0111;
	mem[3576] = 4'b0000;
	mem[3577] = 4'b0000;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b0111;
	mem[3588] = 4'b1100;
	mem[3589] = 4'b1101;
	mem[3590] = 4'b1101;
	mem[3591] = 4'b1101;
	mem[3592] = 4'b1101;
	mem[3593] = 4'b1101;
	mem[3594] = 4'b1101;
	mem[3595] = 4'b1101;
	mem[3596] = 4'b1101;
	mem[3597] = 4'b1101;
	mem[3598] = 4'b1101;
	mem[3599] = 4'b1101;
	mem[3600] = 4'b1101;
	mem[3601] = 4'b1101;
	mem[3602] = 4'b1101;
	mem[3603] = 4'b1101;
	mem[3604] = 4'b1111;
	mem[3605] = 4'b1111;
	mem[3606] = 4'b1111;
	mem[3607] = 4'b1111;
	mem[3608] = 4'b1111;
	mem[3609] = 4'b1111;
	mem[3610] = 4'b1111;
	mem[3611] = 4'b1111;
	mem[3612] = 4'b1111;
	mem[3613] = 4'b1111;
	mem[3614] = 4'b1111;
	mem[3615] = 4'b1111;
	mem[3616] = 4'b1111;
	mem[3617] = 4'b1111;
	mem[3618] = 4'b1111;
	mem[3619] = 4'b1111;
	mem[3620] = 4'b1111;
	mem[3621] = 4'b1000;
	mem[3622] = 4'b0101;
	mem[3623] = 4'b0101;
	mem[3624] = 4'b0101;
	mem[3625] = 4'b0110;
	mem[3626] = 4'b0101;
	mem[3627] = 4'b0101;
	mem[3628] = 4'b0101;
	mem[3629] = 4'b0101;
	mem[3630] = 4'b0101;
	mem[3631] = 4'b0101;
	mem[3632] = 4'b0110;
	mem[3633] = 4'b0110;
	mem[3634] = 4'b0110;
	mem[3635] = 4'b0101;
	mem[3636] = 4'b0101;
	mem[3637] = 4'b0101;
	mem[3638] = 4'b0101;
	mem[3639] = 4'b0110;
	mem[3640] = 4'b0111;
	mem[3641] = 4'b0110;
	mem[3642] = 4'b0110;
	mem[3643] = 4'b0110;
	mem[3644] = 4'b0110;
	mem[3645] = 4'b0110;
	mem[3646] = 4'b0110;
	mem[3647] = 4'b0110;
	mem[3648] = 4'b0110;
	mem[3649] = 4'b0110;
	mem[3650] = 4'b0110;
	mem[3651] = 4'b0110;
	mem[3652] = 4'b0110;
	mem[3653] = 4'b0110;
	mem[3654] = 4'b0110;
	mem[3655] = 4'b1101;
	mem[3656] = 4'b1111;
	mem[3657] = 4'b1111;
	mem[3658] = 4'b1111;
	mem[3659] = 4'b1111;
	mem[3660] = 4'b1111;
	mem[3661] = 4'b1111;
	mem[3662] = 4'b1111;
	mem[3663] = 4'b1111;
	mem[3664] = 4'b1111;
	mem[3665] = 4'b1111;
	mem[3666] = 4'b1111;
	mem[3667] = 4'b1111;
	mem[3668] = 4'b1111;
	mem[3669] = 4'b1111;
	mem[3670] = 4'b1111;
	mem[3671] = 4'b1111;
	mem[3672] = 4'b1111;
	mem[3673] = 4'b1111;
	mem[3674] = 4'b1111;
	mem[3675] = 4'b1110;
	mem[3676] = 4'b1101;
	mem[3677] = 4'b1101;
	mem[3678] = 4'b1110;
	mem[3679] = 4'b1101;
	mem[3680] = 4'b1111;
	mem[3681] = 4'b1111;
	mem[3682] = 4'b1111;
	mem[3683] = 4'b1111;
	mem[3684] = 4'b1111;
	mem[3685] = 4'b1111;
	mem[3686] = 4'b1111;
	mem[3687] = 4'b1110;
	mem[3688] = 4'b1101;
	mem[3689] = 4'b1001;
	mem[3690] = 4'b0110;
	mem[3691] = 4'b0110;
	mem[3692] = 4'b0111;
	mem[3693] = 4'b0111;
	mem[3694] = 4'b0111;
	mem[3695] = 4'b0111;
	mem[3696] = 4'b0111;
	mem[3697] = 4'b0111;
	mem[3698] = 4'b0111;
	mem[3699] = 4'b0111;
	mem[3700] = 4'b0111;
	mem[3701] = 4'b0111;
	mem[3702] = 4'b0111;
	mem[3703] = 4'b0111;
	mem[3704] = 4'b0000;
	mem[3705] = 4'b0000;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b0111;
	mem[3716] = 4'b1100;
	mem[3717] = 4'b1101;
	mem[3718] = 4'b1101;
	mem[3719] = 4'b1101;
	mem[3720] = 4'b1101;
	mem[3721] = 4'b1101;
	mem[3722] = 4'b1101;
	mem[3723] = 4'b1101;
	mem[3724] = 4'b1101;
	mem[3725] = 4'b1101;
	mem[3726] = 4'b1101;
	mem[3727] = 4'b1101;
	mem[3728] = 4'b1101;
	mem[3729] = 4'b1101;
	mem[3730] = 4'b1101;
	mem[3731] = 4'b1101;
	mem[3732] = 4'b1111;
	mem[3733] = 4'b1111;
	mem[3734] = 4'b1111;
	mem[3735] = 4'b1111;
	mem[3736] = 4'b1111;
	mem[3737] = 4'b1111;
	mem[3738] = 4'b1111;
	mem[3739] = 4'b1111;
	mem[3740] = 4'b1111;
	mem[3741] = 4'b1111;
	mem[3742] = 4'b1111;
	mem[3743] = 4'b1111;
	mem[3744] = 4'b1111;
	mem[3745] = 4'b1111;
	mem[3746] = 4'b1111;
	mem[3747] = 4'b1111;
	mem[3748] = 4'b1111;
	mem[3749] = 4'b1000;
	mem[3750] = 4'b0101;
	mem[3751] = 4'b0101;
	mem[3752] = 4'b0101;
	mem[3753] = 4'b0101;
	mem[3754] = 4'b0110;
	mem[3755] = 4'b0101;
	mem[3756] = 4'b0101;
	mem[3757] = 4'b0101;
	mem[3758] = 4'b0110;
	mem[3759] = 4'b0110;
	mem[3760] = 4'b0110;
	mem[3761] = 4'b0110;
	mem[3762] = 4'b0110;
	mem[3763] = 4'b0110;
	mem[3764] = 4'b0101;
	mem[3765] = 4'b0101;
	mem[3766] = 4'b0110;
	mem[3767] = 4'b0111;
	mem[3768] = 4'b0110;
	mem[3769] = 4'b0110;
	mem[3770] = 4'b0110;
	mem[3771] = 4'b0110;
	mem[3772] = 4'b0110;
	mem[3773] = 4'b0110;
	mem[3774] = 4'b0110;
	mem[3775] = 4'b0110;
	mem[3776] = 4'b0110;
	mem[3777] = 4'b0110;
	mem[3778] = 4'b0110;
	mem[3779] = 4'b0110;
	mem[3780] = 4'b0110;
	mem[3781] = 4'b0110;
	mem[3782] = 4'b0110;
	mem[3783] = 4'b1101;
	mem[3784] = 4'b1111;
	mem[3785] = 4'b1111;
	mem[3786] = 4'b1111;
	mem[3787] = 4'b1111;
	mem[3788] = 4'b1111;
	mem[3789] = 4'b1111;
	mem[3790] = 4'b1111;
	mem[3791] = 4'b1111;
	mem[3792] = 4'b1111;
	mem[3793] = 4'b1111;
	mem[3794] = 4'b1111;
	mem[3795] = 4'b1111;
	mem[3796] = 4'b1111;
	mem[3797] = 4'b1111;
	mem[3798] = 4'b1111;
	mem[3799] = 4'b1111;
	mem[3800] = 4'b1111;
	mem[3801] = 4'b1111;
	mem[3802] = 4'b1111;
	mem[3803] = 4'b1101;
	mem[3804] = 4'b1101;
	mem[3805] = 4'b1101;
	mem[3806] = 4'b1101;
	mem[3807] = 4'b1101;
	mem[3808] = 4'b1110;
	mem[3809] = 4'b1111;
	mem[3810] = 4'b1111;
	mem[3811] = 4'b1111;
	mem[3812] = 4'b1111;
	mem[3813] = 4'b1111;
	mem[3814] = 4'b1111;
	mem[3815] = 4'b1111;
	mem[3816] = 4'b1110;
	mem[3817] = 4'b1001;
	mem[3818] = 4'b0110;
	mem[3819] = 4'b0110;
	mem[3820] = 4'b0110;
	mem[3821] = 4'b0111;
	mem[3822] = 4'b0111;
	mem[3823] = 4'b0111;
	mem[3824] = 4'b0111;
	mem[3825] = 4'b0111;
	mem[3826] = 4'b0111;
	mem[3827] = 4'b0111;
	mem[3828] = 4'b0111;
	mem[3829] = 4'b0111;
	mem[3830] = 4'b0111;
	mem[3831] = 4'b0111;
	mem[3832] = 4'b0000;
	mem[3833] = 4'b0000;
	mem[3834] = 4'b0000;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b0111;
	mem[3844] = 4'b1100;
	mem[3845] = 4'b1101;
	mem[3846] = 4'b1101;
	mem[3847] = 4'b1101;
	mem[3848] = 4'b1101;
	mem[3849] = 4'b1101;
	mem[3850] = 4'b1101;
	mem[3851] = 4'b1101;
	mem[3852] = 4'b1101;
	mem[3853] = 4'b1101;
	mem[3854] = 4'b1101;
	mem[3855] = 4'b1101;
	mem[3856] = 4'b1101;
	mem[3857] = 4'b1101;
	mem[3858] = 4'b1101;
	mem[3859] = 4'b1101;
	mem[3860] = 4'b1111;
	mem[3861] = 4'b1111;
	mem[3862] = 4'b1111;
	mem[3863] = 4'b1111;
	mem[3864] = 4'b1111;
	mem[3865] = 4'b1111;
	mem[3866] = 4'b1111;
	mem[3867] = 4'b1111;
	mem[3868] = 4'b1111;
	mem[3869] = 4'b1111;
	mem[3870] = 4'b1111;
	mem[3871] = 4'b1111;
	mem[3872] = 4'b1111;
	mem[3873] = 4'b1111;
	mem[3874] = 4'b1111;
	mem[3875] = 4'b1111;
	mem[3876] = 4'b1111;
	mem[3877] = 4'b1000;
	mem[3878] = 4'b0110;
	mem[3879] = 4'b0101;
	mem[3880] = 4'b0101;
	mem[3881] = 4'b0101;
	mem[3882] = 4'b0101;
	mem[3883] = 4'b0110;
	mem[3884] = 4'b0110;
	mem[3885] = 4'b0110;
	mem[3886] = 4'b0110;
	mem[3887] = 4'b0110;
	mem[3888] = 4'b0110;
	mem[3889] = 4'b0110;
	mem[3890] = 4'b0101;
	mem[3891] = 4'b0110;
	mem[3892] = 4'b0110;
	mem[3893] = 4'b0110;
	mem[3894] = 4'b0111;
	mem[3895] = 4'b0110;
	mem[3896] = 4'b0110;
	mem[3897] = 4'b0110;
	mem[3898] = 4'b0110;
	mem[3899] = 4'b0110;
	mem[3900] = 4'b0110;
	mem[3901] = 4'b0110;
	mem[3902] = 4'b0110;
	mem[3903] = 4'b0110;
	mem[3904] = 4'b0110;
	mem[3905] = 4'b0110;
	mem[3906] = 4'b0110;
	mem[3907] = 4'b0110;
	mem[3908] = 4'b0110;
	mem[3909] = 4'b0110;
	mem[3910] = 4'b0110;
	mem[3911] = 4'b1101;
	mem[3912] = 4'b1111;
	mem[3913] = 4'b1111;
	mem[3914] = 4'b1111;
	mem[3915] = 4'b1111;
	mem[3916] = 4'b1111;
	mem[3917] = 4'b1111;
	mem[3918] = 4'b1111;
	mem[3919] = 4'b1111;
	mem[3920] = 4'b1111;
	mem[3921] = 4'b1111;
	mem[3922] = 4'b1111;
	mem[3923] = 4'b1111;
	mem[3924] = 4'b1111;
	mem[3925] = 4'b1111;
	mem[3926] = 4'b1111;
	mem[3927] = 4'b1111;
	mem[3928] = 4'b1111;
	mem[3929] = 4'b1111;
	mem[3930] = 4'b1111;
	mem[3931] = 4'b1111;
	mem[3932] = 4'b1101;
	mem[3933] = 4'b1101;
	mem[3934] = 4'b1101;
	mem[3935] = 4'b1101;
	mem[3936] = 4'b1101;
	mem[3937] = 4'b1111;
	mem[3938] = 4'b1111;
	mem[3939] = 4'b1111;
	mem[3940] = 4'b1111;
	mem[3941] = 4'b1111;
	mem[3942] = 4'b1111;
	mem[3943] = 4'b1111;
	mem[3944] = 4'b1111;
	mem[3945] = 4'b1001;
	mem[3946] = 4'b0110;
	mem[3947] = 4'b0110;
	mem[3948] = 4'b0110;
	mem[3949] = 4'b0110;
	mem[3950] = 4'b0111;
	mem[3951] = 4'b0111;
	mem[3952] = 4'b0111;
	mem[3953] = 4'b0111;
	mem[3954] = 4'b0111;
	mem[3955] = 4'b0111;
	mem[3956] = 4'b0111;
	mem[3957] = 4'b0111;
	mem[3958] = 4'b0111;
	mem[3959] = 4'b0111;
	mem[3960] = 4'b0000;
	mem[3961] = 4'b0000;
	mem[3962] = 4'b0000;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b0111;
	mem[3972] = 4'b1100;
	mem[3973] = 4'b1101;
	mem[3974] = 4'b1101;
	mem[3975] = 4'b1101;
	mem[3976] = 4'b1101;
	mem[3977] = 4'b1101;
	mem[3978] = 4'b1101;
	mem[3979] = 4'b1101;
	mem[3980] = 4'b1101;
	mem[3981] = 4'b1101;
	mem[3982] = 4'b1101;
	mem[3983] = 4'b1101;
	mem[3984] = 4'b1101;
	mem[3985] = 4'b1101;
	mem[3986] = 4'b1101;
	mem[3987] = 4'b1101;
	mem[3988] = 4'b1111;
	mem[3989] = 4'b1111;
	mem[3990] = 4'b1111;
	mem[3991] = 4'b1111;
	mem[3992] = 4'b1111;
	mem[3993] = 4'b1111;
	mem[3994] = 4'b1111;
	mem[3995] = 4'b1111;
	mem[3996] = 4'b1111;
	mem[3997] = 4'b1111;
	mem[3998] = 4'b1111;
	mem[3999] = 4'b1111;
	mem[4000] = 4'b1111;
	mem[4001] = 4'b1111;
	mem[4002] = 4'b1111;
	mem[4003] = 4'b1111;
	mem[4004] = 4'b1111;
	mem[4005] = 4'b1000;
	mem[4006] = 4'b0101;
	mem[4007] = 4'b0110;
	mem[4008] = 4'b0110;
	mem[4009] = 4'b0101;
	mem[4010] = 4'b0101;
	mem[4011] = 4'b0101;
	mem[4012] = 4'b0110;
	mem[4013] = 4'b0110;
	mem[4014] = 4'b0110;
	mem[4015] = 4'b0110;
	mem[4016] = 4'b0110;
	mem[4017] = 4'b0110;
	mem[4018] = 4'b0101;
	mem[4019] = 4'b0101;
	mem[4020] = 4'b0110;
	mem[4021] = 4'b0110;
	mem[4022] = 4'b0110;
	mem[4023] = 4'b0110;
	mem[4024] = 4'b0110;
	mem[4025] = 4'b0110;
	mem[4026] = 4'b0110;
	mem[4027] = 4'b0110;
	mem[4028] = 4'b0110;
	mem[4029] = 4'b0110;
	mem[4030] = 4'b0110;
	mem[4031] = 4'b0110;
	mem[4032] = 4'b0110;
	mem[4033] = 4'b0110;
	mem[4034] = 4'b0110;
	mem[4035] = 4'b0110;
	mem[4036] = 4'b0110;
	mem[4037] = 4'b0110;
	mem[4038] = 4'b0110;
	mem[4039] = 4'b1101;
	mem[4040] = 4'b1111;
	mem[4041] = 4'b1111;
	mem[4042] = 4'b1111;
	mem[4043] = 4'b1111;
	mem[4044] = 4'b1111;
	mem[4045] = 4'b1111;
	mem[4046] = 4'b1111;
	mem[4047] = 4'b1111;
	mem[4048] = 4'b1111;
	mem[4049] = 4'b1111;
	mem[4050] = 4'b1111;
	mem[4051] = 4'b1111;
	mem[4052] = 4'b1111;
	mem[4053] = 4'b1111;
	mem[4054] = 4'b1111;
	mem[4055] = 4'b1111;
	mem[4056] = 4'b1111;
	mem[4057] = 4'b1111;
	mem[4058] = 4'b1111;
	mem[4059] = 4'b1111;
	mem[4060] = 4'b1111;
	mem[4061] = 4'b1101;
	mem[4062] = 4'b1101;
	mem[4063] = 4'b1101;
	mem[4064] = 4'b1101;
	mem[4065] = 4'b1110;
	mem[4066] = 4'b1111;
	mem[4067] = 4'b1111;
	mem[4068] = 4'b1111;
	mem[4069] = 4'b1111;
	mem[4070] = 4'b1111;
	mem[4071] = 4'b1111;
	mem[4072] = 4'b1111;
	mem[4073] = 4'b1010;
	mem[4074] = 4'b0111;
	mem[4075] = 4'b0110;
	mem[4076] = 4'b0110;
	mem[4077] = 4'b0111;
	mem[4078] = 4'b1000;
	mem[4079] = 4'b0111;
	mem[4080] = 4'b0111;
	mem[4081] = 4'b0111;
	mem[4082] = 4'b0111;
	mem[4083] = 4'b0111;
	mem[4084] = 4'b0111;
	mem[4085] = 4'b0111;
	mem[4086] = 4'b0111;
	mem[4087] = 4'b0111;
	mem[4088] = 4'b0000;
	mem[4089] = 4'b0000;
	mem[4090] = 4'b0000;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_1r (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0111;
	mem[4] = 4'b1100;
	mem[5] = 4'b1101;
	mem[6] = 4'b1101;
	mem[7] = 4'b1101;
	mem[8] = 4'b1101;
	mem[9] = 4'b1101;
	mem[10] = 4'b1101;
	mem[11] = 4'b1101;
	mem[12] = 4'b1101;
	mem[13] = 4'b1101;
	mem[14] = 4'b1101;
	mem[15] = 4'b1101;
	mem[16] = 4'b1101;
	mem[17] = 4'b1101;
	mem[18] = 4'b1101;
	mem[19] = 4'b1101;
	mem[20] = 4'b1111;
	mem[21] = 4'b1111;
	mem[22] = 4'b1111;
	mem[23] = 4'b1111;
	mem[24] = 4'b1111;
	mem[25] = 4'b1111;
	mem[26] = 4'b1111;
	mem[27] = 4'b1111;
	mem[28] = 4'b1111;
	mem[29] = 4'b1111;
	mem[30] = 4'b1111;
	mem[31] = 4'b1111;
	mem[32] = 4'b1111;
	mem[33] = 4'b1111;
	mem[34] = 4'b1111;
	mem[35] = 4'b1111;
	mem[36] = 4'b1111;
	mem[37] = 4'b1000;
	mem[38] = 4'b0101;
	mem[39] = 4'b0101;
	mem[40] = 4'b0110;
	mem[41] = 4'b0110;
	mem[42] = 4'b0101;
	mem[43] = 4'b0101;
	mem[44] = 4'b0110;
	mem[45] = 4'b0110;
	mem[46] = 4'b0110;
	mem[47] = 4'b0110;
	mem[48] = 4'b0110;
	mem[49] = 4'b0101;
	mem[50] = 4'b0101;
	mem[51] = 4'b0110;
	mem[52] = 4'b0110;
	mem[53] = 4'b0110;
	mem[54] = 4'b0110;
	mem[55] = 4'b0110;
	mem[56] = 4'b0110;
	mem[57] = 4'b0110;
	mem[58] = 4'b0110;
	mem[59] = 4'b0110;
	mem[60] = 4'b0110;
	mem[61] = 4'b0110;
	mem[62] = 4'b0110;
	mem[63] = 4'b0110;
	mem[64] = 4'b0110;
	mem[65] = 4'b0110;
	mem[66] = 4'b0110;
	mem[67] = 4'b0110;
	mem[68] = 4'b0110;
	mem[69] = 4'b0110;
	mem[70] = 4'b0110;
	mem[71] = 4'b1101;
	mem[72] = 4'b1111;
	mem[73] = 4'b1111;
	mem[74] = 4'b1111;
	mem[75] = 4'b1111;
	mem[76] = 4'b1111;
	mem[77] = 4'b1111;
	mem[78] = 4'b1111;
	mem[79] = 4'b1111;
	mem[80] = 4'b1111;
	mem[81] = 4'b1111;
	mem[82] = 4'b1111;
	mem[83] = 4'b1111;
	mem[84] = 4'b1111;
	mem[85] = 4'b1111;
	mem[86] = 4'b1111;
	mem[87] = 4'b1111;
	mem[88] = 4'b1111;
	mem[89] = 4'b1111;
	mem[90] = 4'b1111;
	mem[91] = 4'b1111;
	mem[92] = 4'b1111;
	mem[93] = 4'b1111;
	mem[94] = 4'b1101;
	mem[95] = 4'b1101;
	mem[96] = 4'b1101;
	mem[97] = 4'b1101;
	mem[98] = 4'b1110;
	mem[99] = 4'b1111;
	mem[100] = 4'b1111;
	mem[101] = 4'b1111;
	mem[102] = 4'b1111;
	mem[103] = 4'b1111;
	mem[104] = 4'b1111;
	mem[105] = 4'b1010;
	mem[106] = 4'b0111;
	mem[107] = 4'b0111;
	mem[108] = 4'b0111;
	mem[109] = 4'b1000;
	mem[110] = 4'b0111;
	mem[111] = 4'b0111;
	mem[112] = 4'b0111;
	mem[113] = 4'b0111;
	mem[114] = 4'b0111;
	mem[115] = 4'b0111;
	mem[116] = 4'b0111;
	mem[117] = 4'b0111;
	mem[118] = 4'b0111;
	mem[119] = 4'b0111;
	mem[120] = 4'b0000;
	mem[121] = 4'b0000;
	mem[122] = 4'b0000;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b0111;
	mem[132] = 4'b1100;
	mem[133] = 4'b1101;
	mem[134] = 4'b1101;
	mem[135] = 4'b1101;
	mem[136] = 4'b1101;
	mem[137] = 4'b1101;
	mem[138] = 4'b1101;
	mem[139] = 4'b1101;
	mem[140] = 4'b1101;
	mem[141] = 4'b1101;
	mem[142] = 4'b1101;
	mem[143] = 4'b1101;
	mem[144] = 4'b1101;
	mem[145] = 4'b1101;
	mem[146] = 4'b1101;
	mem[147] = 4'b1101;
	mem[148] = 4'b1111;
	mem[149] = 4'b1111;
	mem[150] = 4'b1111;
	mem[151] = 4'b1111;
	mem[152] = 4'b1111;
	mem[153] = 4'b1111;
	mem[154] = 4'b1111;
	mem[155] = 4'b1111;
	mem[156] = 4'b1111;
	mem[157] = 4'b1111;
	mem[158] = 4'b1111;
	mem[159] = 4'b1111;
	mem[160] = 4'b1111;
	mem[161] = 4'b1111;
	mem[162] = 4'b1111;
	mem[163] = 4'b1111;
	mem[164] = 4'b1111;
	mem[165] = 4'b1000;
	mem[166] = 4'b0110;
	mem[167] = 4'b0110;
	mem[168] = 4'b0110;
	mem[169] = 4'b0110;
	mem[170] = 4'b0110;
	mem[171] = 4'b0101;
	mem[172] = 4'b0101;
	mem[173] = 4'b0110;
	mem[174] = 4'b0110;
	mem[175] = 4'b0110;
	mem[176] = 4'b0101;
	mem[177] = 4'b0101;
	mem[178] = 4'b0110;
	mem[179] = 4'b0111;
	mem[180] = 4'b0110;
	mem[181] = 4'b0110;
	mem[182] = 4'b0110;
	mem[183] = 4'b0110;
	mem[184] = 4'b0110;
	mem[185] = 4'b0110;
	mem[186] = 4'b0110;
	mem[187] = 4'b0110;
	mem[188] = 4'b0110;
	mem[189] = 4'b0110;
	mem[190] = 4'b0110;
	mem[191] = 4'b0110;
	mem[192] = 4'b0110;
	mem[193] = 4'b0110;
	mem[194] = 4'b0110;
	mem[195] = 4'b0110;
	mem[196] = 4'b0110;
	mem[197] = 4'b0110;
	mem[198] = 4'b0110;
	mem[199] = 4'b1101;
	mem[200] = 4'b1111;
	mem[201] = 4'b1111;
	mem[202] = 4'b1111;
	mem[203] = 4'b1111;
	mem[204] = 4'b1111;
	mem[205] = 4'b1111;
	mem[206] = 4'b1111;
	mem[207] = 4'b1111;
	mem[208] = 4'b1111;
	mem[209] = 4'b1111;
	mem[210] = 4'b1111;
	mem[211] = 4'b1111;
	mem[212] = 4'b1111;
	mem[213] = 4'b1111;
	mem[214] = 4'b1110;
	mem[215] = 4'b1110;
	mem[216] = 4'b1111;
	mem[217] = 4'b1111;
	mem[218] = 4'b1111;
	mem[219] = 4'b1111;
	mem[220] = 4'b1111;
	mem[221] = 4'b1111;
	mem[222] = 4'b1111;
	mem[223] = 4'b1101;
	mem[224] = 4'b1101;
	mem[225] = 4'b1101;
	mem[226] = 4'b1101;
	mem[227] = 4'b1110;
	mem[228] = 4'b1111;
	mem[229] = 4'b1111;
	mem[230] = 4'b1111;
	mem[231] = 4'b1111;
	mem[232] = 4'b1111;
	mem[233] = 4'b1010;
	mem[234] = 4'b0111;
	mem[235] = 4'b0111;
	mem[236] = 4'b1000;
	mem[237] = 4'b0111;
	mem[238] = 4'b0111;
	mem[239] = 4'b0111;
	mem[240] = 4'b0111;
	mem[241] = 4'b0111;
	mem[242] = 4'b0111;
	mem[243] = 4'b0111;
	mem[244] = 4'b0111;
	mem[245] = 4'b0111;
	mem[246] = 4'b0111;
	mem[247] = 4'b0111;
	mem[248] = 4'b0000;
	mem[249] = 4'b0000;
	mem[250] = 4'b0000;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0111;
	mem[260] = 4'b1100;
	mem[261] = 4'b1101;
	mem[262] = 4'b1101;
	mem[263] = 4'b1101;
	mem[264] = 4'b1101;
	mem[265] = 4'b1101;
	mem[266] = 4'b1101;
	mem[267] = 4'b1101;
	mem[268] = 4'b1101;
	mem[269] = 4'b1101;
	mem[270] = 4'b1101;
	mem[271] = 4'b1101;
	mem[272] = 4'b1101;
	mem[273] = 4'b1101;
	mem[274] = 4'b1101;
	mem[275] = 4'b1101;
	mem[276] = 4'b1111;
	mem[277] = 4'b1111;
	mem[278] = 4'b1111;
	mem[279] = 4'b1111;
	mem[280] = 4'b1111;
	mem[281] = 4'b1111;
	mem[282] = 4'b1111;
	mem[283] = 4'b1111;
	mem[284] = 4'b1111;
	mem[285] = 4'b1111;
	mem[286] = 4'b1111;
	mem[287] = 4'b1111;
	mem[288] = 4'b1111;
	mem[289] = 4'b1111;
	mem[290] = 4'b1111;
	mem[291] = 4'b1111;
	mem[292] = 4'b1111;
	mem[293] = 4'b1000;
	mem[294] = 4'b0110;
	mem[295] = 4'b0110;
	mem[296] = 4'b0110;
	mem[297] = 4'b0110;
	mem[298] = 4'b0110;
	mem[299] = 4'b0110;
	mem[300] = 4'b0101;
	mem[301] = 4'b0101;
	mem[302] = 4'b0110;
	mem[303] = 4'b0101;
	mem[304] = 4'b0101;
	mem[305] = 4'b0110;
	mem[306] = 4'b0111;
	mem[307] = 4'b0110;
	mem[308] = 4'b0110;
	mem[309] = 4'b0110;
	mem[310] = 4'b0110;
	mem[311] = 4'b0110;
	mem[312] = 4'b0110;
	mem[313] = 4'b0110;
	mem[314] = 4'b0110;
	mem[315] = 4'b0110;
	mem[316] = 4'b0110;
	mem[317] = 4'b0110;
	mem[318] = 4'b0110;
	mem[319] = 4'b0110;
	mem[320] = 4'b0110;
	mem[321] = 4'b0110;
	mem[322] = 4'b0110;
	mem[323] = 4'b0110;
	mem[324] = 4'b0110;
	mem[325] = 4'b0110;
	mem[326] = 4'b0110;
	mem[327] = 4'b1101;
	mem[328] = 4'b1111;
	mem[329] = 4'b1111;
	mem[330] = 4'b1111;
	mem[331] = 4'b1111;
	mem[332] = 4'b1111;
	mem[333] = 4'b1111;
	mem[334] = 4'b1111;
	mem[335] = 4'b1111;
	mem[336] = 4'b1111;
	mem[337] = 4'b1111;
	mem[338] = 4'b1111;
	mem[339] = 4'b1111;
	mem[340] = 4'b1110;
	mem[341] = 4'b1101;
	mem[342] = 4'b1101;
	mem[343] = 4'b1101;
	mem[344] = 4'b1101;
	mem[345] = 4'b1110;
	mem[346] = 4'b1111;
	mem[347] = 4'b1111;
	mem[348] = 4'b1111;
	mem[349] = 4'b1111;
	mem[350] = 4'b1111;
	mem[351] = 4'b1111;
	mem[352] = 4'b1101;
	mem[353] = 4'b1101;
	mem[354] = 4'b1101;
	mem[355] = 4'b1101;
	mem[356] = 4'b1110;
	mem[357] = 4'b1111;
	mem[358] = 4'b1111;
	mem[359] = 4'b1111;
	mem[360] = 4'b1111;
	mem[361] = 4'b1010;
	mem[362] = 4'b0111;
	mem[363] = 4'b0111;
	mem[364] = 4'b0111;
	mem[365] = 4'b0111;
	mem[366] = 4'b0111;
	mem[367] = 4'b0111;
	mem[368] = 4'b0111;
	mem[369] = 4'b0111;
	mem[370] = 4'b0111;
	mem[371] = 4'b0111;
	mem[372] = 4'b0111;
	mem[373] = 4'b0111;
	mem[374] = 4'b0111;
	mem[375] = 4'b0111;
	mem[376] = 4'b0000;
	mem[377] = 4'b0000;
	mem[378] = 4'b0000;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0111;
	mem[388] = 4'b1100;
	mem[389] = 4'b1101;
	mem[390] = 4'b1101;
	mem[391] = 4'b1101;
	mem[392] = 4'b1101;
	mem[393] = 4'b1101;
	mem[394] = 4'b1101;
	mem[395] = 4'b1101;
	mem[396] = 4'b1101;
	mem[397] = 4'b1101;
	mem[398] = 4'b1101;
	mem[399] = 4'b1101;
	mem[400] = 4'b1101;
	mem[401] = 4'b1101;
	mem[402] = 4'b1101;
	mem[403] = 4'b1101;
	mem[404] = 4'b1111;
	mem[405] = 4'b1111;
	mem[406] = 4'b1111;
	mem[407] = 4'b1111;
	mem[408] = 4'b1111;
	mem[409] = 4'b1111;
	mem[410] = 4'b1111;
	mem[411] = 4'b1111;
	mem[412] = 4'b1111;
	mem[413] = 4'b1111;
	mem[414] = 4'b1111;
	mem[415] = 4'b1111;
	mem[416] = 4'b1111;
	mem[417] = 4'b1111;
	mem[418] = 4'b1111;
	mem[419] = 4'b1111;
	mem[420] = 4'b1111;
	mem[421] = 4'b1000;
	mem[422] = 4'b0110;
	mem[423] = 4'b0110;
	mem[424] = 4'b0101;
	mem[425] = 4'b0101;
	mem[426] = 4'b0110;
	mem[427] = 4'b0110;
	mem[428] = 4'b0110;
	mem[429] = 4'b0101;
	mem[430] = 4'b0101;
	mem[431] = 4'b0101;
	mem[432] = 4'b0110;
	mem[433] = 4'b0111;
	mem[434] = 4'b0110;
	mem[435] = 4'b0110;
	mem[436] = 4'b0110;
	mem[437] = 4'b0110;
	mem[438] = 4'b0110;
	mem[439] = 4'b0110;
	mem[440] = 4'b0110;
	mem[441] = 4'b0110;
	mem[442] = 4'b0110;
	mem[443] = 4'b0110;
	mem[444] = 4'b0110;
	mem[445] = 4'b0110;
	mem[446] = 4'b0110;
	mem[447] = 4'b0110;
	mem[448] = 4'b0110;
	mem[449] = 4'b0110;
	mem[450] = 4'b0110;
	mem[451] = 4'b0110;
	mem[452] = 4'b0110;
	mem[453] = 4'b0110;
	mem[454] = 4'b0110;
	mem[455] = 4'b1101;
	mem[456] = 4'b1111;
	mem[457] = 4'b1111;
	mem[458] = 4'b1111;
	mem[459] = 4'b1111;
	mem[460] = 4'b1111;
	mem[461] = 4'b1111;
	mem[462] = 4'b1111;
	mem[463] = 4'b1111;
	mem[464] = 4'b1111;
	mem[465] = 4'b1111;
	mem[466] = 4'b1111;
	mem[467] = 4'b1110;
	mem[468] = 4'b1101;
	mem[469] = 4'b1101;
	mem[470] = 4'b1101;
	mem[471] = 4'b1101;
	mem[472] = 4'b1101;
	mem[473] = 4'b1101;
	mem[474] = 4'b1101;
	mem[475] = 4'b1111;
	mem[476] = 4'b1111;
	mem[477] = 4'b1111;
	mem[478] = 4'b1111;
	mem[479] = 4'b1111;
	mem[480] = 4'b1111;
	mem[481] = 4'b1101;
	mem[482] = 4'b1101;
	mem[483] = 4'b1101;
	mem[484] = 4'b1101;
	mem[485] = 4'b1110;
	mem[486] = 4'b1111;
	mem[487] = 4'b1111;
	mem[488] = 4'b1111;
	mem[489] = 4'b1010;
	mem[490] = 4'b0111;
	mem[491] = 4'b0111;
	mem[492] = 4'b0111;
	mem[493] = 4'b0111;
	mem[494] = 4'b0111;
	mem[495] = 4'b0111;
	mem[496] = 4'b0111;
	mem[497] = 4'b0111;
	mem[498] = 4'b0111;
	mem[499] = 4'b0111;
	mem[500] = 4'b0111;
	mem[501] = 4'b0111;
	mem[502] = 4'b0111;
	mem[503] = 4'b0111;
	mem[504] = 4'b0000;
	mem[505] = 4'b0000;
	mem[506] = 4'b0000;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0111;
	mem[516] = 4'b1100;
	mem[517] = 4'b1101;
	mem[518] = 4'b1101;
	mem[519] = 4'b1101;
	mem[520] = 4'b1101;
	mem[521] = 4'b1101;
	mem[522] = 4'b1101;
	mem[523] = 4'b1101;
	mem[524] = 4'b1101;
	mem[525] = 4'b1101;
	mem[526] = 4'b1101;
	mem[527] = 4'b1101;
	mem[528] = 4'b1101;
	mem[529] = 4'b1101;
	mem[530] = 4'b1101;
	mem[531] = 4'b1101;
	mem[532] = 4'b1111;
	mem[533] = 4'b1111;
	mem[534] = 4'b1111;
	mem[535] = 4'b1111;
	mem[536] = 4'b1111;
	mem[537] = 4'b1111;
	mem[538] = 4'b1111;
	mem[539] = 4'b1111;
	mem[540] = 4'b1111;
	mem[541] = 4'b1111;
	mem[542] = 4'b1111;
	mem[543] = 4'b1111;
	mem[544] = 4'b1111;
	mem[545] = 4'b1111;
	mem[546] = 4'b1111;
	mem[547] = 4'b1111;
	mem[548] = 4'b1111;
	mem[549] = 4'b1000;
	mem[550] = 4'b0110;
	mem[551] = 4'b0101;
	mem[552] = 4'b0101;
	mem[553] = 4'b0101;
	mem[554] = 4'b0110;
	mem[555] = 4'b0110;
	mem[556] = 4'b0110;
	mem[557] = 4'b0110;
	mem[558] = 4'b0101;
	mem[559] = 4'b0110;
	mem[560] = 4'b0111;
	mem[561] = 4'b0110;
	mem[562] = 4'b0110;
	mem[563] = 4'b0110;
	mem[564] = 4'b0110;
	mem[565] = 4'b0110;
	mem[566] = 4'b0110;
	mem[567] = 4'b0110;
	mem[568] = 4'b0110;
	mem[569] = 4'b0110;
	mem[570] = 4'b0110;
	mem[571] = 4'b0110;
	mem[572] = 4'b0110;
	mem[573] = 4'b0110;
	mem[574] = 4'b0110;
	mem[575] = 4'b0110;
	mem[576] = 4'b0110;
	mem[577] = 4'b0110;
	mem[578] = 4'b0110;
	mem[579] = 4'b0110;
	mem[580] = 4'b0110;
	mem[581] = 4'b0110;
	mem[582] = 4'b0110;
	mem[583] = 4'b1101;
	mem[584] = 4'b1111;
	mem[585] = 4'b1111;
	mem[586] = 4'b1111;
	mem[587] = 4'b1111;
	mem[588] = 4'b1111;
	mem[589] = 4'b1111;
	mem[590] = 4'b1111;
	mem[591] = 4'b1111;
	mem[592] = 4'b1111;
	mem[593] = 4'b1111;
	mem[594] = 4'b1110;
	mem[595] = 4'b1101;
	mem[596] = 4'b1101;
	mem[597] = 4'b1101;
	mem[598] = 4'b1101;
	mem[599] = 4'b1101;
	mem[600] = 4'b1101;
	mem[601] = 4'b1101;
	mem[602] = 4'b1101;
	mem[603] = 4'b1101;
	mem[604] = 4'b1111;
	mem[605] = 4'b1111;
	mem[606] = 4'b1111;
	mem[607] = 4'b1111;
	mem[608] = 4'b1111;
	mem[609] = 4'b1111;
	mem[610] = 4'b1101;
	mem[611] = 4'b1101;
	mem[612] = 4'b1101;
	mem[613] = 4'b1101;
	mem[614] = 4'b1110;
	mem[615] = 4'b1111;
	mem[616] = 4'b1111;
	mem[617] = 4'b1010;
	mem[618] = 4'b0111;
	mem[619] = 4'b0111;
	mem[620] = 4'b0111;
	mem[621] = 4'b0111;
	mem[622] = 4'b0111;
	mem[623] = 4'b0111;
	mem[624] = 4'b0111;
	mem[625] = 4'b0111;
	mem[626] = 4'b0111;
	mem[627] = 4'b0111;
	mem[628] = 4'b0111;
	mem[629] = 4'b0111;
	mem[630] = 4'b0111;
	mem[631] = 4'b0111;
	mem[632] = 4'b0000;
	mem[633] = 4'b0000;
	mem[634] = 4'b0000;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0111;
	mem[644] = 4'b1100;
	mem[645] = 4'b1101;
	mem[646] = 4'b1101;
	mem[647] = 4'b1101;
	mem[648] = 4'b1101;
	mem[649] = 4'b1101;
	mem[650] = 4'b1101;
	mem[651] = 4'b1101;
	mem[652] = 4'b1101;
	mem[653] = 4'b1101;
	mem[654] = 4'b1101;
	mem[655] = 4'b1101;
	mem[656] = 4'b1101;
	mem[657] = 4'b1101;
	mem[658] = 4'b1101;
	mem[659] = 4'b1101;
	mem[660] = 4'b1111;
	mem[661] = 4'b1111;
	mem[662] = 4'b1111;
	mem[663] = 4'b1111;
	mem[664] = 4'b1111;
	mem[665] = 4'b1111;
	mem[666] = 4'b1111;
	mem[667] = 4'b1111;
	mem[668] = 4'b1111;
	mem[669] = 4'b1111;
	mem[670] = 4'b1111;
	mem[671] = 4'b1111;
	mem[672] = 4'b1111;
	mem[673] = 4'b1111;
	mem[674] = 4'b1111;
	mem[675] = 4'b1111;
	mem[676] = 4'b1111;
	mem[677] = 4'b1000;
	mem[678] = 4'b0101;
	mem[679] = 4'b0101;
	mem[680] = 4'b0101;
	mem[681] = 4'b0110;
	mem[682] = 4'b0111;
	mem[683] = 4'b0110;
	mem[684] = 4'b0110;
	mem[685] = 4'b0110;
	mem[686] = 4'b0110;
	mem[687] = 4'b0111;
	mem[688] = 4'b0110;
	mem[689] = 4'b0110;
	mem[690] = 4'b0110;
	mem[691] = 4'b0110;
	mem[692] = 4'b0110;
	mem[693] = 4'b0110;
	mem[694] = 4'b0110;
	mem[695] = 4'b0110;
	mem[696] = 4'b0110;
	mem[697] = 4'b0110;
	mem[698] = 4'b0110;
	mem[699] = 4'b0110;
	mem[700] = 4'b0110;
	mem[701] = 4'b0110;
	mem[702] = 4'b0110;
	mem[703] = 4'b0110;
	mem[704] = 4'b0110;
	mem[705] = 4'b0110;
	mem[706] = 4'b0110;
	mem[707] = 4'b0110;
	mem[708] = 4'b0110;
	mem[709] = 4'b0110;
	mem[710] = 4'b0110;
	mem[711] = 4'b1101;
	mem[712] = 4'b1111;
	mem[713] = 4'b1111;
	mem[714] = 4'b1111;
	mem[715] = 4'b1111;
	mem[716] = 4'b1111;
	mem[717] = 4'b1111;
	mem[718] = 4'b1111;
	mem[719] = 4'b1111;
	mem[720] = 4'b1111;
	mem[721] = 4'b1110;
	mem[722] = 4'b1101;
	mem[723] = 4'b1101;
	mem[724] = 4'b1101;
	mem[725] = 4'b1110;
	mem[726] = 4'b1111;
	mem[727] = 4'b1111;
	mem[728] = 4'b1110;
	mem[729] = 4'b1101;
	mem[730] = 4'b1101;
	mem[731] = 4'b1101;
	mem[732] = 4'b1101;
	mem[733] = 4'b1111;
	mem[734] = 4'b1111;
	mem[735] = 4'b1111;
	mem[736] = 4'b1111;
	mem[737] = 4'b1111;
	mem[738] = 4'b1111;
	mem[739] = 4'b1101;
	mem[740] = 4'b1101;
	mem[741] = 4'b1101;
	mem[742] = 4'b1101;
	mem[743] = 4'b1111;
	mem[744] = 4'b1111;
	mem[745] = 4'b1010;
	mem[746] = 4'b0111;
	mem[747] = 4'b0111;
	mem[748] = 4'b0111;
	mem[749] = 4'b0111;
	mem[750] = 4'b0111;
	mem[751] = 4'b0111;
	mem[752] = 4'b0111;
	mem[753] = 4'b0111;
	mem[754] = 4'b0111;
	mem[755] = 4'b0111;
	mem[756] = 4'b0111;
	mem[757] = 4'b0111;
	mem[758] = 4'b1000;
	mem[759] = 4'b1000;
	mem[760] = 4'b0000;
	mem[761] = 4'b0000;
	mem[762] = 4'b0000;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0111;
	mem[772] = 4'b1100;
	mem[773] = 4'b1101;
	mem[774] = 4'b1101;
	mem[775] = 4'b1101;
	mem[776] = 4'b1101;
	mem[777] = 4'b1101;
	mem[778] = 4'b1101;
	mem[779] = 4'b1101;
	mem[780] = 4'b1101;
	mem[781] = 4'b1101;
	mem[782] = 4'b1101;
	mem[783] = 4'b1101;
	mem[784] = 4'b1101;
	mem[785] = 4'b1101;
	mem[786] = 4'b1101;
	mem[787] = 4'b1101;
	mem[788] = 4'b1111;
	mem[789] = 4'b1111;
	mem[790] = 4'b1111;
	mem[791] = 4'b1111;
	mem[792] = 4'b1111;
	mem[793] = 4'b1111;
	mem[794] = 4'b1111;
	mem[795] = 4'b1111;
	mem[796] = 4'b1111;
	mem[797] = 4'b1111;
	mem[798] = 4'b1111;
	mem[799] = 4'b1111;
	mem[800] = 4'b1111;
	mem[801] = 4'b1110;
	mem[802] = 4'b1110;
	mem[803] = 4'b1110;
	mem[804] = 4'b1111;
	mem[805] = 4'b1000;
	mem[806] = 4'b0110;
	mem[807] = 4'b0101;
	mem[808] = 4'b0110;
	mem[809] = 4'b0111;
	mem[810] = 4'b0110;
	mem[811] = 4'b0110;
	mem[812] = 4'b0110;
	mem[813] = 4'b0110;
	mem[814] = 4'b0110;
	mem[815] = 4'b0110;
	mem[816] = 4'b0110;
	mem[817] = 4'b0110;
	mem[818] = 4'b0110;
	mem[819] = 4'b0110;
	mem[820] = 4'b0110;
	mem[821] = 4'b0110;
	mem[822] = 4'b0110;
	mem[823] = 4'b0110;
	mem[824] = 4'b0110;
	mem[825] = 4'b0110;
	mem[826] = 4'b0110;
	mem[827] = 4'b0110;
	mem[828] = 4'b0110;
	mem[829] = 4'b0110;
	mem[830] = 4'b0110;
	mem[831] = 4'b0110;
	mem[832] = 4'b0110;
	mem[833] = 4'b0110;
	mem[834] = 4'b0110;
	mem[835] = 4'b0110;
	mem[836] = 4'b0110;
	mem[837] = 4'b0110;
	mem[838] = 4'b0110;
	mem[839] = 4'b1101;
	mem[840] = 4'b1111;
	mem[841] = 4'b1111;
	mem[842] = 4'b1111;
	mem[843] = 4'b1111;
	mem[844] = 4'b1111;
	mem[845] = 4'b1111;
	mem[846] = 4'b1111;
	mem[847] = 4'b1111;
	mem[848] = 4'b1111;
	mem[849] = 4'b1101;
	mem[850] = 4'b1101;
	mem[851] = 4'b1101;
	mem[852] = 4'b1110;
	mem[853] = 4'b1111;
	mem[854] = 4'b1111;
	mem[855] = 4'b1111;
	mem[856] = 4'b1110;
	mem[857] = 4'b1101;
	mem[858] = 4'b1101;
	mem[859] = 4'b1101;
	mem[860] = 4'b1101;
	mem[861] = 4'b1101;
	mem[862] = 4'b1111;
	mem[863] = 4'b1111;
	mem[864] = 4'b1111;
	mem[865] = 4'b1111;
	mem[866] = 4'b1111;
	mem[867] = 4'b1111;
	mem[868] = 4'b1101;
	mem[869] = 4'b1101;
	mem[870] = 4'b1110;
	mem[871] = 4'b1111;
	mem[872] = 4'b1111;
	mem[873] = 4'b1010;
	mem[874] = 4'b0111;
	mem[875] = 4'b0111;
	mem[876] = 4'b0111;
	mem[877] = 4'b0111;
	mem[878] = 4'b0110;
	mem[879] = 4'b0101;
	mem[880] = 4'b0100;
	mem[881] = 4'b0100;
	mem[882] = 4'b0011;
	mem[883] = 4'b0010;
	mem[884] = 4'b0010;
	mem[885] = 4'b0001;
	mem[886] = 4'b0000;
	mem[887] = 4'b0000;
	mem[888] = 4'b0000;
	mem[889] = 4'b0000;
	mem[890] = 4'b0000;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0111;
	mem[900] = 4'b1100;
	mem[901] = 4'b1101;
	mem[902] = 4'b1101;
	mem[903] = 4'b1101;
	mem[904] = 4'b1101;
	mem[905] = 4'b1101;
	mem[906] = 4'b1101;
	mem[907] = 4'b1101;
	mem[908] = 4'b1101;
	mem[909] = 4'b1101;
	mem[910] = 4'b1101;
	mem[911] = 4'b1101;
	mem[912] = 4'b1101;
	mem[913] = 4'b1101;
	mem[914] = 4'b1101;
	mem[915] = 4'b1101;
	mem[916] = 4'b1111;
	mem[917] = 4'b1111;
	mem[918] = 4'b1111;
	mem[919] = 4'b1111;
	mem[920] = 4'b1111;
	mem[921] = 4'b1111;
	mem[922] = 4'b1111;
	mem[923] = 4'b1111;
	mem[924] = 4'b1111;
	mem[925] = 4'b1111;
	mem[926] = 4'b1111;
	mem[927] = 4'b1111;
	mem[928] = 4'b1110;
	mem[929] = 4'b1101;
	mem[930] = 4'b1101;
	mem[931] = 4'b1111;
	mem[932] = 4'b1111;
	mem[933] = 4'b1000;
	mem[934] = 4'b0110;
	mem[935] = 4'b0110;
	mem[936] = 4'b0111;
	mem[937] = 4'b0110;
	mem[938] = 4'b0110;
	mem[939] = 4'b0110;
	mem[940] = 4'b0110;
	mem[941] = 4'b0110;
	mem[942] = 4'b0110;
	mem[943] = 4'b0110;
	mem[944] = 4'b0110;
	mem[945] = 4'b0110;
	mem[946] = 4'b0110;
	mem[947] = 4'b0110;
	mem[948] = 4'b0110;
	mem[949] = 4'b0110;
	mem[950] = 4'b0110;
	mem[951] = 4'b0110;
	mem[952] = 4'b0110;
	mem[953] = 4'b0110;
	mem[954] = 4'b0110;
	mem[955] = 4'b0110;
	mem[956] = 4'b0110;
	mem[957] = 4'b0110;
	mem[958] = 4'b0110;
	mem[959] = 4'b0110;
	mem[960] = 4'b0110;
	mem[961] = 4'b0110;
	mem[962] = 4'b0110;
	mem[963] = 4'b0110;
	mem[964] = 4'b0110;
	mem[965] = 4'b0110;
	mem[966] = 4'b0110;
	mem[967] = 4'b1101;
	mem[968] = 4'b1111;
	mem[969] = 4'b1111;
	mem[970] = 4'b1111;
	mem[971] = 4'b1111;
	mem[972] = 4'b1111;
	mem[973] = 4'b1111;
	mem[974] = 4'b1111;
	mem[975] = 4'b1111;
	mem[976] = 4'b1110;
	mem[977] = 4'b1101;
	mem[978] = 4'b1101;
	mem[979] = 4'b1110;
	mem[980] = 4'b1111;
	mem[981] = 4'b1111;
	mem[982] = 4'b1111;
	mem[983] = 4'b1111;
	mem[984] = 4'b1101;
	mem[985] = 4'b1101;
	mem[986] = 4'b1101;
	mem[987] = 4'b1101;
	mem[988] = 4'b1101;
	mem[989] = 4'b1101;
	mem[990] = 4'b1101;
	mem[991] = 4'b1111;
	mem[992] = 4'b1111;
	mem[993] = 4'b1111;
	mem[994] = 4'b1111;
	mem[995] = 4'b1111;
	mem[996] = 4'b1111;
	mem[997] = 4'b1110;
	mem[998] = 4'b1111;
	mem[999] = 4'b1111;
	mem[1000] = 4'b1111;
	mem[1001] = 4'b1000;
	mem[1002] = 4'b0010;
	mem[1003] = 4'b0001;
	mem[1004] = 4'b0000;
	mem[1005] = 4'b0000;
	mem[1006] = 4'b0000;
	mem[1007] = 4'b0000;
	mem[1008] = 4'b0000;
	mem[1009] = 4'b0000;
	mem[1010] = 4'b0000;
	mem[1011] = 4'b0000;
	mem[1012] = 4'b0000;
	mem[1013] = 4'b0000;
	mem[1014] = 4'b0000;
	mem[1015] = 4'b0000;
	mem[1016] = 4'b0000;
	mem[1017] = 4'b0000;
	mem[1018] = 4'b0000;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0111;
	mem[1028] = 4'b1100;
	mem[1029] = 4'b1101;
	mem[1030] = 4'b1101;
	mem[1031] = 4'b1101;
	mem[1032] = 4'b1101;
	mem[1033] = 4'b1101;
	mem[1034] = 4'b1101;
	mem[1035] = 4'b1101;
	mem[1036] = 4'b1101;
	mem[1037] = 4'b1101;
	mem[1038] = 4'b1101;
	mem[1039] = 4'b1101;
	mem[1040] = 4'b1101;
	mem[1041] = 4'b1101;
	mem[1042] = 4'b1101;
	mem[1043] = 4'b1101;
	mem[1044] = 4'b1111;
	mem[1045] = 4'b1111;
	mem[1046] = 4'b1111;
	mem[1047] = 4'b1111;
	mem[1048] = 4'b1111;
	mem[1049] = 4'b1111;
	mem[1050] = 4'b1111;
	mem[1051] = 4'b1111;
	mem[1052] = 4'b1111;
	mem[1053] = 4'b1111;
	mem[1054] = 4'b1111;
	mem[1055] = 4'b1110;
	mem[1056] = 4'b1101;
	mem[1057] = 4'b1111;
	mem[1058] = 4'b1111;
	mem[1059] = 4'b1111;
	mem[1060] = 4'b1111;
	mem[1061] = 4'b1000;
	mem[1062] = 4'b0110;
	mem[1063] = 4'b0110;
	mem[1064] = 4'b0110;
	mem[1065] = 4'b0110;
	mem[1066] = 4'b0110;
	mem[1067] = 4'b0110;
	mem[1068] = 4'b0110;
	mem[1069] = 4'b0110;
	mem[1070] = 4'b0110;
	mem[1071] = 4'b0110;
	mem[1072] = 4'b0110;
	mem[1073] = 4'b0110;
	mem[1074] = 4'b0110;
	mem[1075] = 4'b0110;
	mem[1076] = 4'b0110;
	mem[1077] = 4'b0110;
	mem[1078] = 4'b0110;
	mem[1079] = 4'b0110;
	mem[1080] = 4'b0110;
	mem[1081] = 4'b0110;
	mem[1082] = 4'b0110;
	mem[1083] = 4'b0110;
	mem[1084] = 4'b0110;
	mem[1085] = 4'b0110;
	mem[1086] = 4'b0110;
	mem[1087] = 4'b0110;
	mem[1088] = 4'b0110;
	mem[1089] = 4'b0110;
	mem[1090] = 4'b0110;
	mem[1091] = 4'b0110;
	mem[1092] = 4'b0110;
	mem[1093] = 4'b0111;
	mem[1094] = 4'b0111;
	mem[1095] = 4'b1101;
	mem[1096] = 4'b1111;
	mem[1097] = 4'b1111;
	mem[1098] = 4'b1111;
	mem[1099] = 4'b1111;
	mem[1100] = 4'b1111;
	mem[1101] = 4'b1111;
	mem[1102] = 4'b1111;
	mem[1103] = 4'b1111;
	mem[1104] = 4'b1110;
	mem[1105] = 4'b1101;
	mem[1106] = 4'b1101;
	mem[1107] = 4'b1110;
	mem[1108] = 4'b1111;
	mem[1109] = 4'b1111;
	mem[1110] = 4'b1111;
	mem[1111] = 4'b1110;
	mem[1112] = 4'b1101;
	mem[1113] = 4'b1110;
	mem[1114] = 4'b1111;
	mem[1115] = 4'b1101;
	mem[1116] = 4'b1101;
	mem[1117] = 4'b1101;
	mem[1118] = 4'b1101;
	mem[1119] = 4'b1101;
	mem[1120] = 4'b1111;
	mem[1121] = 4'b1111;
	mem[1122] = 4'b1111;
	mem[1123] = 4'b1111;
	mem[1124] = 4'b1111;
	mem[1125] = 4'b1111;
	mem[1126] = 4'b1111;
	mem[1127] = 4'b1111;
	mem[1128] = 4'b1111;
	mem[1129] = 4'b0110;
	mem[1130] = 4'b0000;
	mem[1131] = 4'b0000;
	mem[1132] = 4'b0000;
	mem[1133] = 4'b0000;
	mem[1134] = 4'b0000;
	mem[1135] = 4'b0000;
	mem[1136] = 4'b0000;
	mem[1137] = 4'b0000;
	mem[1138] = 4'b0000;
	mem[1139] = 4'b0000;
	mem[1140] = 4'b0000;
	mem[1141] = 4'b0000;
	mem[1142] = 4'b0000;
	mem[1143] = 4'b0000;
	mem[1144] = 4'b0000;
	mem[1145] = 4'b0000;
	mem[1146] = 4'b0000;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0111;
	mem[1156] = 4'b1100;
	mem[1157] = 4'b1101;
	mem[1158] = 4'b1101;
	mem[1159] = 4'b1101;
	mem[1160] = 4'b1101;
	mem[1161] = 4'b1101;
	mem[1162] = 4'b1101;
	mem[1163] = 4'b1101;
	mem[1164] = 4'b1101;
	mem[1165] = 4'b1101;
	mem[1166] = 4'b1101;
	mem[1167] = 4'b1101;
	mem[1168] = 4'b1101;
	mem[1169] = 4'b1101;
	mem[1170] = 4'b1101;
	mem[1171] = 4'b1101;
	mem[1172] = 4'b1111;
	mem[1173] = 4'b1111;
	mem[1174] = 4'b1111;
	mem[1175] = 4'b1111;
	mem[1176] = 4'b1111;
	mem[1177] = 4'b1111;
	mem[1178] = 4'b1111;
	mem[1179] = 4'b1111;
	mem[1180] = 4'b1111;
	mem[1181] = 4'b1111;
	mem[1182] = 4'b1110;
	mem[1183] = 4'b1101;
	mem[1184] = 4'b1111;
	mem[1185] = 4'b1111;
	mem[1186] = 4'b1111;
	mem[1187] = 4'b1110;
	mem[1188] = 4'b1101;
	mem[1189] = 4'b0111;
	mem[1190] = 4'b0101;
	mem[1191] = 4'b0110;
	mem[1192] = 4'b0110;
	mem[1193] = 4'b0110;
	mem[1194] = 4'b0110;
	mem[1195] = 4'b0110;
	mem[1196] = 4'b0110;
	mem[1197] = 4'b0110;
	mem[1198] = 4'b0110;
	mem[1199] = 4'b0110;
	mem[1200] = 4'b0110;
	mem[1201] = 4'b0110;
	mem[1202] = 4'b0110;
	mem[1203] = 4'b0110;
	mem[1204] = 4'b0110;
	mem[1205] = 4'b0110;
	mem[1206] = 4'b0110;
	mem[1207] = 4'b0110;
	mem[1208] = 4'b0110;
	mem[1209] = 4'b0110;
	mem[1210] = 4'b0110;
	mem[1211] = 4'b0110;
	mem[1212] = 4'b0110;
	mem[1213] = 4'b0110;
	mem[1214] = 4'b0110;
	mem[1215] = 4'b0110;
	mem[1216] = 4'b0110;
	mem[1217] = 4'b0110;
	mem[1218] = 4'b0110;
	mem[1219] = 4'b0111;
	mem[1220] = 4'b0111;
	mem[1221] = 4'b0111;
	mem[1222] = 4'b0111;
	mem[1223] = 4'b1101;
	mem[1224] = 4'b1111;
	mem[1225] = 4'b1111;
	mem[1226] = 4'b1111;
	mem[1227] = 4'b1111;
	mem[1228] = 4'b1111;
	mem[1229] = 4'b1111;
	mem[1230] = 4'b1111;
	mem[1231] = 4'b1111;
	mem[1232] = 4'b1110;
	mem[1233] = 4'b1101;
	mem[1234] = 4'b1101;
	mem[1235] = 4'b1110;
	mem[1236] = 4'b1111;
	mem[1237] = 4'b1111;
	mem[1238] = 4'b1110;
	mem[1239] = 4'b1101;
	mem[1240] = 4'b1101;
	mem[1241] = 4'b1111;
	mem[1242] = 4'b1111;
	mem[1243] = 4'b1111;
	mem[1244] = 4'b1101;
	mem[1245] = 4'b1101;
	mem[1246] = 4'b1101;
	mem[1247] = 4'b1101;
	mem[1248] = 4'b1101;
	mem[1249] = 4'b1110;
	mem[1250] = 4'b1111;
	mem[1251] = 4'b1111;
	mem[1252] = 4'b1111;
	mem[1253] = 4'b1111;
	mem[1254] = 4'b1111;
	mem[1255] = 4'b1111;
	mem[1256] = 4'b1111;
	mem[1257] = 4'b0110;
	mem[1258] = 4'b0000;
	mem[1259] = 4'b0000;
	mem[1260] = 4'b0000;
	mem[1261] = 4'b0000;
	mem[1262] = 4'b0000;
	mem[1263] = 4'b0000;
	mem[1264] = 4'b0000;
	mem[1265] = 4'b0000;
	mem[1266] = 4'b0000;
	mem[1267] = 4'b0000;
	mem[1268] = 4'b0000;
	mem[1269] = 4'b0000;
	mem[1270] = 4'b0000;
	mem[1271] = 4'b0000;
	mem[1272] = 4'b0000;
	mem[1273] = 4'b0000;
	mem[1274] = 4'b0000;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0111;
	mem[1284] = 4'b1100;
	mem[1285] = 4'b1101;
	mem[1286] = 4'b1101;
	mem[1287] = 4'b1101;
	mem[1288] = 4'b1101;
	mem[1289] = 4'b1101;
	mem[1290] = 4'b1101;
	mem[1291] = 4'b1101;
	mem[1292] = 4'b1101;
	mem[1293] = 4'b1101;
	mem[1294] = 4'b1101;
	mem[1295] = 4'b1101;
	mem[1296] = 4'b1101;
	mem[1297] = 4'b1101;
	mem[1298] = 4'b1101;
	mem[1299] = 4'b1101;
	mem[1300] = 4'b1111;
	mem[1301] = 4'b1111;
	mem[1302] = 4'b1111;
	mem[1303] = 4'b1111;
	mem[1304] = 4'b1111;
	mem[1305] = 4'b1111;
	mem[1306] = 4'b1111;
	mem[1307] = 4'b1111;
	mem[1308] = 4'b1111;
	mem[1309] = 4'b1111;
	mem[1310] = 4'b1110;
	mem[1311] = 4'b1101;
	mem[1312] = 4'b1110;
	mem[1313] = 4'b1110;
	mem[1314] = 4'b1101;
	mem[1315] = 4'b1101;
	mem[1316] = 4'b1110;
	mem[1317] = 4'b1000;
	mem[1318] = 4'b0101;
	mem[1319] = 4'b0110;
	mem[1320] = 4'b0110;
	mem[1321] = 4'b0110;
	mem[1322] = 4'b0110;
	mem[1323] = 4'b0110;
	mem[1324] = 4'b0110;
	mem[1325] = 4'b0110;
	mem[1326] = 4'b0110;
	mem[1327] = 4'b0110;
	mem[1328] = 4'b0110;
	mem[1329] = 4'b0110;
	mem[1330] = 4'b0110;
	mem[1331] = 4'b0110;
	mem[1332] = 4'b0110;
	mem[1333] = 4'b0110;
	mem[1334] = 4'b0110;
	mem[1335] = 4'b0110;
	mem[1336] = 4'b0110;
	mem[1337] = 4'b0110;
	mem[1338] = 4'b0110;
	mem[1339] = 4'b0110;
	mem[1340] = 4'b0110;
	mem[1341] = 4'b0110;
	mem[1342] = 4'b0110;
	mem[1343] = 4'b0110;
	mem[1344] = 4'b0110;
	mem[1345] = 4'b0111;
	mem[1346] = 4'b0111;
	mem[1347] = 4'b0111;
	mem[1348] = 4'b0111;
	mem[1349] = 4'b0111;
	mem[1350] = 4'b0111;
	mem[1351] = 4'b1101;
	mem[1352] = 4'b1111;
	mem[1353] = 4'b1111;
	mem[1354] = 4'b1111;
	mem[1355] = 4'b1111;
	mem[1356] = 4'b1111;
	mem[1357] = 4'b1111;
	mem[1358] = 4'b1111;
	mem[1359] = 4'b1111;
	mem[1360] = 4'b1111;
	mem[1361] = 4'b1101;
	mem[1362] = 4'b1110;
	mem[1363] = 4'b1111;
	mem[1364] = 4'b1111;
	mem[1365] = 4'b1111;
	mem[1366] = 4'b1101;
	mem[1367] = 4'b1101;
	mem[1368] = 4'b1110;
	mem[1369] = 4'b1111;
	mem[1370] = 4'b1111;
	mem[1371] = 4'b1111;
	mem[1372] = 4'b1110;
	mem[1373] = 4'b1101;
	mem[1374] = 4'b1101;
	mem[1375] = 4'b1101;
	mem[1376] = 4'b1101;
	mem[1377] = 4'b1101;
	mem[1378] = 4'b1111;
	mem[1379] = 4'b1111;
	mem[1380] = 4'b1111;
	mem[1381] = 4'b1111;
	mem[1382] = 4'b1111;
	mem[1383] = 4'b1111;
	mem[1384] = 4'b1111;
	mem[1385] = 4'b0110;
	mem[1386] = 4'b0000;
	mem[1387] = 4'b0000;
	mem[1388] = 4'b0000;
	mem[1389] = 4'b0000;
	mem[1390] = 4'b0000;
	mem[1391] = 4'b0000;
	mem[1392] = 4'b0000;
	mem[1393] = 4'b0000;
	mem[1394] = 4'b0000;
	mem[1395] = 4'b0000;
	mem[1396] = 4'b0000;
	mem[1397] = 4'b0000;
	mem[1398] = 4'b0000;
	mem[1399] = 4'b0000;
	mem[1400] = 4'b0000;
	mem[1401] = 4'b0000;
	mem[1402] = 4'b0000;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0111;
	mem[1412] = 4'b1100;
	mem[1413] = 4'b1101;
	mem[1414] = 4'b1101;
	mem[1415] = 4'b1101;
	mem[1416] = 4'b1101;
	mem[1417] = 4'b1101;
	mem[1418] = 4'b1101;
	mem[1419] = 4'b1101;
	mem[1420] = 4'b1101;
	mem[1421] = 4'b1101;
	mem[1422] = 4'b1101;
	mem[1423] = 4'b1101;
	mem[1424] = 4'b1101;
	mem[1425] = 4'b1101;
	mem[1426] = 4'b1101;
	mem[1427] = 4'b1101;
	mem[1428] = 4'b1111;
	mem[1429] = 4'b1111;
	mem[1430] = 4'b1111;
	mem[1431] = 4'b1111;
	mem[1432] = 4'b1111;
	mem[1433] = 4'b1111;
	mem[1434] = 4'b1111;
	mem[1435] = 4'b1111;
	mem[1436] = 4'b1111;
	mem[1437] = 4'b1111;
	mem[1438] = 4'b1111;
	mem[1439] = 4'b1101;
	mem[1440] = 4'b1101;
	mem[1441] = 4'b1101;
	mem[1442] = 4'b1101;
	mem[1443] = 4'b1110;
	mem[1444] = 4'b1111;
	mem[1445] = 4'b1001;
	mem[1446] = 4'b0101;
	mem[1447] = 4'b0110;
	mem[1448] = 4'b0111;
	mem[1449] = 4'b0110;
	mem[1450] = 4'b0110;
	mem[1451] = 4'b0110;
	mem[1452] = 4'b0110;
	mem[1453] = 4'b0110;
	mem[1454] = 4'b0110;
	mem[1455] = 4'b0110;
	mem[1456] = 4'b0110;
	mem[1457] = 4'b0110;
	mem[1458] = 4'b0110;
	mem[1459] = 4'b0110;
	mem[1460] = 4'b0110;
	mem[1461] = 4'b0110;
	mem[1462] = 4'b0110;
	mem[1463] = 4'b0110;
	mem[1464] = 4'b0110;
	mem[1465] = 4'b0110;
	mem[1466] = 4'b0110;
	mem[1467] = 4'b0110;
	mem[1468] = 4'b0110;
	mem[1469] = 4'b0110;
	mem[1470] = 4'b0110;
	mem[1471] = 4'b0111;
	mem[1472] = 4'b0111;
	mem[1473] = 4'b0111;
	mem[1474] = 4'b0111;
	mem[1475] = 4'b0111;
	mem[1476] = 4'b0111;
	mem[1477] = 4'b0111;
	mem[1478] = 4'b0111;
	mem[1479] = 4'b1101;
	mem[1480] = 4'b1111;
	mem[1481] = 4'b1111;
	mem[1482] = 4'b1111;
	mem[1483] = 4'b1111;
	mem[1484] = 4'b1111;
	mem[1485] = 4'b1111;
	mem[1486] = 4'b1111;
	mem[1487] = 4'b1111;
	mem[1488] = 4'b1111;
	mem[1489] = 4'b1111;
	mem[1490] = 4'b1111;
	mem[1491] = 4'b1111;
	mem[1492] = 4'b1111;
	mem[1493] = 4'b1110;
	mem[1494] = 4'b1101;
	mem[1495] = 4'b1101;
	mem[1496] = 4'b1111;
	mem[1497] = 4'b1111;
	mem[1498] = 4'b1111;
	mem[1499] = 4'b1111;
	mem[1500] = 4'b1110;
	mem[1501] = 4'b1101;
	mem[1502] = 4'b1110;
	mem[1503] = 4'b1101;
	mem[1504] = 4'b1110;
	mem[1505] = 4'b1111;
	mem[1506] = 4'b1111;
	mem[1507] = 4'b1111;
	mem[1508] = 4'b1111;
	mem[1509] = 4'b1111;
	mem[1510] = 4'b1111;
	mem[1511] = 4'b1111;
	mem[1512] = 4'b1111;
	mem[1513] = 4'b0110;
	mem[1514] = 4'b0000;
	mem[1515] = 4'b0000;
	mem[1516] = 4'b0000;
	mem[1517] = 4'b0000;
	mem[1518] = 4'b0000;
	mem[1519] = 4'b0000;
	mem[1520] = 4'b0000;
	mem[1521] = 4'b0000;
	mem[1522] = 4'b0000;
	mem[1523] = 4'b0000;
	mem[1524] = 4'b0000;
	mem[1525] = 4'b0000;
	mem[1526] = 4'b0000;
	mem[1527] = 4'b0000;
	mem[1528] = 4'b0000;
	mem[1529] = 4'b0000;
	mem[1530] = 4'b0000;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0111;
	mem[1540] = 4'b1100;
	mem[1541] = 4'b1101;
	mem[1542] = 4'b1101;
	mem[1543] = 4'b1101;
	mem[1544] = 4'b1101;
	mem[1545] = 4'b1101;
	mem[1546] = 4'b1101;
	mem[1547] = 4'b1101;
	mem[1548] = 4'b1101;
	mem[1549] = 4'b1101;
	mem[1550] = 4'b1101;
	mem[1551] = 4'b1101;
	mem[1552] = 4'b1101;
	mem[1553] = 4'b1101;
	mem[1554] = 4'b1101;
	mem[1555] = 4'b1101;
	mem[1556] = 4'b1111;
	mem[1557] = 4'b1111;
	mem[1558] = 4'b1111;
	mem[1559] = 4'b1111;
	mem[1560] = 4'b1111;
	mem[1561] = 4'b1111;
	mem[1562] = 4'b1111;
	mem[1563] = 4'b1111;
	mem[1564] = 4'b1111;
	mem[1565] = 4'b1111;
	mem[1566] = 4'b1111;
	mem[1567] = 4'b1111;
	mem[1568] = 4'b1110;
	mem[1569] = 4'b1110;
	mem[1570] = 4'b1111;
	mem[1571] = 4'b1111;
	mem[1572] = 4'b1111;
	mem[1573] = 4'b1000;
	mem[1574] = 4'b0101;
	mem[1575] = 4'b0111;
	mem[1576] = 4'b0110;
	mem[1577] = 4'b0110;
	mem[1578] = 4'b0110;
	mem[1579] = 4'b0110;
	mem[1580] = 4'b0110;
	mem[1581] = 4'b0110;
	mem[1582] = 4'b0110;
	mem[1583] = 4'b0110;
	mem[1584] = 4'b0110;
	mem[1585] = 4'b0110;
	mem[1586] = 4'b0110;
	mem[1587] = 4'b0110;
	mem[1588] = 4'b0110;
	mem[1589] = 4'b0110;
	mem[1590] = 4'b0110;
	mem[1591] = 4'b0110;
	mem[1592] = 4'b0110;
	mem[1593] = 4'b0110;
	mem[1594] = 4'b0110;
	mem[1595] = 4'b0110;
	mem[1596] = 4'b0110;
	mem[1597] = 4'b0111;
	mem[1598] = 4'b0111;
	mem[1599] = 4'b0111;
	mem[1600] = 4'b0111;
	mem[1601] = 4'b0111;
	mem[1602] = 4'b0111;
	mem[1603] = 4'b0111;
	mem[1604] = 4'b0111;
	mem[1605] = 4'b0111;
	mem[1606] = 4'b0111;
	mem[1607] = 4'b1101;
	mem[1608] = 4'b1111;
	mem[1609] = 4'b1111;
	mem[1610] = 4'b1111;
	mem[1611] = 4'b1111;
	mem[1612] = 4'b1111;
	mem[1613] = 4'b1111;
	mem[1614] = 4'b1111;
	mem[1615] = 4'b1111;
	mem[1616] = 4'b1111;
	mem[1617] = 4'b1111;
	mem[1618] = 4'b1111;
	mem[1619] = 4'b1111;
	mem[1620] = 4'b1111;
	mem[1621] = 4'b1101;
	mem[1622] = 4'b1101;
	mem[1623] = 4'b1110;
	mem[1624] = 4'b1111;
	mem[1625] = 4'b1111;
	mem[1626] = 4'b1111;
	mem[1627] = 4'b1111;
	mem[1628] = 4'b1110;
	mem[1629] = 4'b1101;
	mem[1630] = 4'b1111;
	mem[1631] = 4'b1111;
	mem[1632] = 4'b1111;
	mem[1633] = 4'b1111;
	mem[1634] = 4'b1111;
	mem[1635] = 4'b1111;
	mem[1636] = 4'b1111;
	mem[1637] = 4'b1111;
	mem[1638] = 4'b1111;
	mem[1639] = 4'b1111;
	mem[1640] = 4'b1111;
	mem[1641] = 4'b0110;
	mem[1642] = 4'b0000;
	mem[1643] = 4'b0000;
	mem[1644] = 4'b0000;
	mem[1645] = 4'b0000;
	mem[1646] = 4'b0000;
	mem[1647] = 4'b0000;
	mem[1648] = 4'b0000;
	mem[1649] = 4'b0000;
	mem[1650] = 4'b0000;
	mem[1651] = 4'b0000;
	mem[1652] = 4'b0000;
	mem[1653] = 4'b0000;
	mem[1654] = 4'b0000;
	mem[1655] = 4'b0000;
	mem[1656] = 4'b0000;
	mem[1657] = 4'b0000;
	mem[1658] = 4'b0000;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0111;
	mem[1668] = 4'b1100;
	mem[1669] = 4'b1101;
	mem[1670] = 4'b1101;
	mem[1671] = 4'b1101;
	mem[1672] = 4'b1101;
	mem[1673] = 4'b1101;
	mem[1674] = 4'b1101;
	mem[1675] = 4'b1101;
	mem[1676] = 4'b1101;
	mem[1677] = 4'b1101;
	mem[1678] = 4'b1101;
	mem[1679] = 4'b1101;
	mem[1680] = 4'b1101;
	mem[1681] = 4'b1101;
	mem[1682] = 4'b1101;
	mem[1683] = 4'b1101;
	mem[1684] = 4'b1111;
	mem[1685] = 4'b1111;
	mem[1686] = 4'b1111;
	mem[1687] = 4'b1111;
	mem[1688] = 4'b1111;
	mem[1689] = 4'b1111;
	mem[1690] = 4'b1110;
	mem[1691] = 4'b1101;
	mem[1692] = 4'b1101;
	mem[1693] = 4'b1111;
	mem[1694] = 4'b1111;
	mem[1695] = 4'b1111;
	mem[1696] = 4'b1111;
	mem[1697] = 4'b1111;
	mem[1698] = 4'b1111;
	mem[1699] = 4'b1110;
	mem[1700] = 4'b1110;
	mem[1701] = 4'b0111;
	mem[1702] = 4'b0110;
	mem[1703] = 4'b0111;
	mem[1704] = 4'b0110;
	mem[1705] = 4'b0110;
	mem[1706] = 4'b0110;
	mem[1707] = 4'b0110;
	mem[1708] = 4'b0110;
	mem[1709] = 4'b0110;
	mem[1710] = 4'b0110;
	mem[1711] = 4'b0110;
	mem[1712] = 4'b0110;
	mem[1713] = 4'b0110;
	mem[1714] = 4'b0110;
	mem[1715] = 4'b0110;
	mem[1716] = 4'b0110;
	mem[1717] = 4'b0110;
	mem[1718] = 4'b0110;
	mem[1719] = 4'b0110;
	mem[1720] = 4'b0110;
	mem[1721] = 4'b0110;
	mem[1722] = 4'b0110;
	mem[1723] = 4'b0110;
	mem[1724] = 4'b0111;
	mem[1725] = 4'b0111;
	mem[1726] = 4'b0111;
	mem[1727] = 4'b0111;
	mem[1728] = 4'b0111;
	mem[1729] = 4'b0111;
	mem[1730] = 4'b0111;
	mem[1731] = 4'b0111;
	mem[1732] = 4'b0111;
	mem[1733] = 4'b0111;
	mem[1734] = 4'b0111;
	mem[1735] = 4'b1101;
	mem[1736] = 4'b1111;
	mem[1737] = 4'b1111;
	mem[1738] = 4'b1111;
	mem[1739] = 4'b1111;
	mem[1740] = 4'b1111;
	mem[1741] = 4'b1111;
	mem[1742] = 4'b1111;
	mem[1743] = 4'b1111;
	mem[1744] = 4'b1111;
	mem[1745] = 4'b1111;
	mem[1746] = 4'b1111;
	mem[1747] = 4'b1111;
	mem[1748] = 4'b1110;
	mem[1749] = 4'b1101;
	mem[1750] = 4'b1101;
	mem[1751] = 4'b1101;
	mem[1752] = 4'b1111;
	mem[1753] = 4'b1111;
	mem[1754] = 4'b1111;
	mem[1755] = 4'b1110;
	mem[1756] = 4'b1101;
	mem[1757] = 4'b1101;
	mem[1758] = 4'b1111;
	mem[1759] = 4'b1111;
	mem[1760] = 4'b1111;
	mem[1761] = 4'b1111;
	mem[1762] = 4'b1111;
	mem[1763] = 4'b1111;
	mem[1764] = 4'b1111;
	mem[1765] = 4'b1111;
	mem[1766] = 4'b1111;
	mem[1767] = 4'b1111;
	mem[1768] = 4'b1111;
	mem[1769] = 4'b0110;
	mem[1770] = 4'b0000;
	mem[1771] = 4'b0000;
	mem[1772] = 4'b0000;
	mem[1773] = 4'b0000;
	mem[1774] = 4'b0000;
	mem[1775] = 4'b0000;
	mem[1776] = 4'b0000;
	mem[1777] = 4'b0000;
	mem[1778] = 4'b0000;
	mem[1779] = 4'b0000;
	mem[1780] = 4'b0000;
	mem[1781] = 4'b0000;
	mem[1782] = 4'b0000;
	mem[1783] = 4'b0000;
	mem[1784] = 4'b0000;
	mem[1785] = 4'b0000;
	mem[1786] = 4'b0000;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0111;
	mem[1796] = 4'b1100;
	mem[1797] = 4'b1101;
	mem[1798] = 4'b1101;
	mem[1799] = 4'b1101;
	mem[1800] = 4'b1101;
	mem[1801] = 4'b1101;
	mem[1802] = 4'b1101;
	mem[1803] = 4'b1101;
	mem[1804] = 4'b1101;
	mem[1805] = 4'b1101;
	mem[1806] = 4'b1101;
	mem[1807] = 4'b1101;
	mem[1808] = 4'b1101;
	mem[1809] = 4'b1101;
	mem[1810] = 4'b1101;
	mem[1811] = 4'b1101;
	mem[1812] = 4'b1111;
	mem[1813] = 4'b1111;
	mem[1814] = 4'b1111;
	mem[1815] = 4'b1111;
	mem[1816] = 4'b1111;
	mem[1817] = 4'b1110;
	mem[1818] = 4'b1101;
	mem[1819] = 4'b1101;
	mem[1820] = 4'b1101;
	mem[1821] = 4'b1101;
	mem[1822] = 4'b1110;
	mem[1823] = 4'b1111;
	mem[1824] = 4'b1111;
	mem[1825] = 4'b1111;
	mem[1826] = 4'b1101;
	mem[1827] = 4'b1101;
	mem[1828] = 4'b1101;
	mem[1829] = 4'b1000;
	mem[1830] = 4'b0111;
	mem[1831] = 4'b0110;
	mem[1832] = 4'b0110;
	mem[1833] = 4'b0110;
	mem[1834] = 4'b0110;
	mem[1835] = 4'b0110;
	mem[1836] = 4'b0110;
	mem[1837] = 4'b0110;
	mem[1838] = 4'b0110;
	mem[1839] = 4'b0110;
	mem[1840] = 4'b0110;
	mem[1841] = 4'b0110;
	mem[1842] = 4'b0110;
	mem[1843] = 4'b0110;
	mem[1844] = 4'b0110;
	mem[1845] = 4'b0110;
	mem[1846] = 4'b0110;
	mem[1847] = 4'b0110;
	mem[1848] = 4'b0110;
	mem[1849] = 4'b0110;
	mem[1850] = 4'b0111;
	mem[1851] = 4'b0111;
	mem[1852] = 4'b0111;
	mem[1853] = 4'b0111;
	mem[1854] = 4'b0111;
	mem[1855] = 4'b0111;
	mem[1856] = 4'b0111;
	mem[1857] = 4'b0111;
	mem[1858] = 4'b0111;
	mem[1859] = 4'b0111;
	mem[1860] = 4'b0111;
	mem[1861] = 4'b0101;
	mem[1862] = 4'b0011;
	mem[1863] = 4'b1100;
	mem[1864] = 4'b1111;
	mem[1865] = 4'b1111;
	mem[1866] = 4'b1111;
	mem[1867] = 4'b1111;
	mem[1868] = 4'b1111;
	mem[1869] = 4'b1111;
	mem[1870] = 4'b1111;
	mem[1871] = 4'b1111;
	mem[1872] = 4'b1111;
	mem[1873] = 4'b1111;
	mem[1874] = 4'b1111;
	mem[1875] = 4'b1111;
	mem[1876] = 4'b1111;
	mem[1877] = 4'b1101;
	mem[1878] = 4'b1101;
	mem[1879] = 4'b1101;
	mem[1880] = 4'b1110;
	mem[1881] = 4'b1110;
	mem[1882] = 4'b1110;
	mem[1883] = 4'b1101;
	mem[1884] = 4'b1101;
	mem[1885] = 4'b1110;
	mem[1886] = 4'b1111;
	mem[1887] = 4'b1111;
	mem[1888] = 4'b1111;
	mem[1889] = 4'b1111;
	mem[1890] = 4'b1111;
	mem[1891] = 4'b1111;
	mem[1892] = 4'b1111;
	mem[1893] = 4'b1111;
	mem[1894] = 4'b1111;
	mem[1895] = 4'b1111;
	mem[1896] = 4'b1111;
	mem[1897] = 4'b0110;
	mem[1898] = 4'b0000;
	mem[1899] = 4'b0000;
	mem[1900] = 4'b0000;
	mem[1901] = 4'b0000;
	mem[1902] = 4'b0000;
	mem[1903] = 4'b0000;
	mem[1904] = 4'b0000;
	mem[1905] = 4'b0000;
	mem[1906] = 4'b0000;
	mem[1907] = 4'b0000;
	mem[1908] = 4'b0000;
	mem[1909] = 4'b0000;
	mem[1910] = 4'b0000;
	mem[1911] = 4'b0000;
	mem[1912] = 4'b0000;
	mem[1913] = 4'b0000;
	mem[1914] = 4'b0000;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0111;
	mem[1924] = 4'b1100;
	mem[1925] = 4'b1101;
	mem[1926] = 4'b1101;
	mem[1927] = 4'b1101;
	mem[1928] = 4'b1101;
	mem[1929] = 4'b1101;
	mem[1930] = 4'b1101;
	mem[1931] = 4'b1101;
	mem[1932] = 4'b1101;
	mem[1933] = 4'b1101;
	mem[1934] = 4'b1101;
	mem[1935] = 4'b1101;
	mem[1936] = 4'b1101;
	mem[1937] = 4'b1101;
	mem[1938] = 4'b1101;
	mem[1939] = 4'b1110;
	mem[1940] = 4'b1111;
	mem[1941] = 4'b1111;
	mem[1942] = 4'b1111;
	mem[1943] = 4'b1111;
	mem[1944] = 4'b1111;
	mem[1945] = 4'b1101;
	mem[1946] = 4'b1110;
	mem[1947] = 4'b1111;
	mem[1948] = 4'b1110;
	mem[1949] = 4'b1101;
	mem[1950] = 4'b1101;
	mem[1951] = 4'b1110;
	mem[1952] = 4'b1111;
	mem[1953] = 4'b1111;
	mem[1954] = 4'b1111;
	mem[1955] = 4'b1111;
	mem[1956] = 4'b1111;
	mem[1957] = 4'b1001;
	mem[1958] = 4'b0110;
	mem[1959] = 4'b0110;
	mem[1960] = 4'b0110;
	mem[1961] = 4'b0110;
	mem[1962] = 4'b0110;
	mem[1963] = 4'b0110;
	mem[1964] = 4'b0110;
	mem[1965] = 4'b0110;
	mem[1966] = 4'b0110;
	mem[1967] = 4'b0110;
	mem[1968] = 4'b0110;
	mem[1969] = 4'b0110;
	mem[1970] = 4'b0110;
	mem[1971] = 4'b0110;
	mem[1972] = 4'b0110;
	mem[1973] = 4'b0110;
	mem[1974] = 4'b0110;
	mem[1975] = 4'b0110;
	mem[1976] = 4'b0111;
	mem[1977] = 4'b0111;
	mem[1978] = 4'b0111;
	mem[1979] = 4'b0111;
	mem[1980] = 4'b0111;
	mem[1981] = 4'b0111;
	mem[1982] = 4'b0111;
	mem[1983] = 4'b0111;
	mem[1984] = 4'b0110;
	mem[1985] = 4'b0110;
	mem[1986] = 4'b0100;
	mem[1987] = 4'b0010;
	mem[1988] = 4'b0000;
	mem[1989] = 4'b0000;
	mem[1990] = 4'b0000;
	mem[1991] = 4'b1100;
	mem[1992] = 4'b1111;
	mem[1993] = 4'b1111;
	mem[1994] = 4'b1111;
	mem[1995] = 4'b1111;
	mem[1996] = 4'b1111;
	mem[1997] = 4'b1111;
	mem[1998] = 4'b1111;
	mem[1999] = 4'b1111;
	mem[2000] = 4'b1111;
	mem[2001] = 4'b1111;
	mem[2002] = 4'b1111;
	mem[2003] = 4'b1111;
	mem[2004] = 4'b1111;
	mem[2005] = 4'b1101;
	mem[2006] = 4'b1101;
	mem[2007] = 4'b1101;
	mem[2008] = 4'b1101;
	mem[2009] = 4'b1101;
	mem[2010] = 4'b1101;
	mem[2011] = 4'b1101;
	mem[2012] = 4'b1101;
	mem[2013] = 4'b1111;
	mem[2014] = 4'b1111;
	mem[2015] = 4'b1111;
	mem[2016] = 4'b1111;
	mem[2017] = 4'b1111;
	mem[2018] = 4'b1111;
	mem[2019] = 4'b1111;
	mem[2020] = 4'b1111;
	mem[2021] = 4'b1111;
	mem[2022] = 4'b1111;
	mem[2023] = 4'b1111;
	mem[2024] = 4'b1111;
	mem[2025] = 4'b0110;
	mem[2026] = 4'b0000;
	mem[2027] = 4'b0000;
	mem[2028] = 4'b0000;
	mem[2029] = 4'b0000;
	mem[2030] = 4'b0000;
	mem[2031] = 4'b0000;
	mem[2032] = 4'b0000;
	mem[2033] = 4'b0000;
	mem[2034] = 4'b0000;
	mem[2035] = 4'b0000;
	mem[2036] = 4'b0000;
	mem[2037] = 4'b0000;
	mem[2038] = 4'b0000;
	mem[2039] = 4'b0000;
	mem[2040] = 4'b0000;
	mem[2041] = 4'b0000;
	mem[2042] = 4'b0000;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0111;
	mem[2052] = 4'b1100;
	mem[2053] = 4'b1101;
	mem[2054] = 4'b1101;
	mem[2055] = 4'b1101;
	mem[2056] = 4'b1101;
	mem[2057] = 4'b1101;
	mem[2058] = 4'b1101;
	mem[2059] = 4'b1101;
	mem[2060] = 4'b1101;
	mem[2061] = 4'b1101;
	mem[2062] = 4'b1101;
	mem[2063] = 4'b1101;
	mem[2064] = 4'b1101;
	mem[2065] = 4'b1101;
	mem[2066] = 4'b1110;
	mem[2067] = 4'b1110;
	mem[2068] = 4'b1111;
	mem[2069] = 4'b1111;
	mem[2070] = 4'b1111;
	mem[2071] = 4'b1110;
	mem[2072] = 4'b1110;
	mem[2073] = 4'b1110;
	mem[2074] = 4'b1111;
	mem[2075] = 4'b1111;
	mem[2076] = 4'b1111;
	mem[2077] = 4'b1111;
	mem[2078] = 4'b1101;
	mem[2079] = 4'b1101;
	mem[2080] = 4'b1110;
	mem[2081] = 4'b1111;
	mem[2082] = 4'b1111;
	mem[2083] = 4'b1111;
	mem[2084] = 4'b1111;
	mem[2085] = 4'b1000;
	mem[2086] = 4'b0110;
	mem[2087] = 4'b0110;
	mem[2088] = 4'b0110;
	mem[2089] = 4'b0110;
	mem[2090] = 4'b0110;
	mem[2091] = 4'b0110;
	mem[2092] = 4'b0110;
	mem[2093] = 4'b0110;
	mem[2094] = 4'b0110;
	mem[2095] = 4'b0110;
	mem[2096] = 4'b0110;
	mem[2097] = 4'b0110;
	mem[2098] = 4'b0110;
	mem[2099] = 4'b0110;
	mem[2100] = 4'b0110;
	mem[2101] = 4'b0110;
	mem[2102] = 4'b0111;
	mem[2103] = 4'b0111;
	mem[2104] = 4'b0111;
	mem[2105] = 4'b0111;
	mem[2106] = 4'b0111;
	mem[2107] = 4'b0111;
	mem[2108] = 4'b0111;
	mem[2109] = 4'b0111;
	mem[2110] = 4'b0110;
	mem[2111] = 4'b0011;
	mem[2112] = 4'b0001;
	mem[2113] = 4'b0000;
	mem[2114] = 4'b0000;
	mem[2115] = 4'b0000;
	mem[2116] = 4'b0000;
	mem[2117] = 4'b0000;
	mem[2118] = 4'b0000;
	mem[2119] = 4'b1100;
	mem[2120] = 4'b1111;
	mem[2121] = 4'b1111;
	mem[2122] = 4'b1111;
	mem[2123] = 4'b1111;
	mem[2124] = 4'b1111;
	mem[2125] = 4'b1111;
	mem[2126] = 4'b1111;
	mem[2127] = 4'b1111;
	mem[2128] = 4'b1111;
	mem[2129] = 4'b1111;
	mem[2130] = 4'b1111;
	mem[2131] = 4'b1111;
	mem[2132] = 4'b1111;
	mem[2133] = 4'b1111;
	mem[2134] = 4'b1101;
	mem[2135] = 4'b1101;
	mem[2136] = 4'b1101;
	mem[2137] = 4'b1101;
	mem[2138] = 4'b1101;
	mem[2139] = 4'b1101;
	mem[2140] = 4'b1111;
	mem[2141] = 4'b1111;
	mem[2142] = 4'b1111;
	mem[2143] = 4'b1111;
	mem[2144] = 4'b1111;
	mem[2145] = 4'b1111;
	mem[2146] = 4'b1111;
	mem[2147] = 4'b1111;
	mem[2148] = 4'b1111;
	mem[2149] = 4'b1111;
	mem[2150] = 4'b1111;
	mem[2151] = 4'b1111;
	mem[2152] = 4'b1111;
	mem[2153] = 4'b0110;
	mem[2154] = 4'b0000;
	mem[2155] = 4'b0000;
	mem[2156] = 4'b0000;
	mem[2157] = 4'b0000;
	mem[2158] = 4'b0000;
	mem[2159] = 4'b0000;
	mem[2160] = 4'b0000;
	mem[2161] = 4'b0000;
	mem[2162] = 4'b0000;
	mem[2163] = 4'b0000;
	mem[2164] = 4'b0000;
	mem[2165] = 4'b0000;
	mem[2166] = 4'b0000;
	mem[2167] = 4'b0000;
	mem[2168] = 4'b0000;
	mem[2169] = 4'b0000;
	mem[2170] = 4'b0000;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0111;
	mem[2180] = 4'b1100;
	mem[2181] = 4'b1101;
	mem[2182] = 4'b1101;
	mem[2183] = 4'b1101;
	mem[2184] = 4'b1101;
	mem[2185] = 4'b1101;
	mem[2186] = 4'b1101;
	mem[2187] = 4'b1101;
	mem[2188] = 4'b1101;
	mem[2189] = 4'b1101;
	mem[2190] = 4'b1101;
	mem[2191] = 4'b1101;
	mem[2192] = 4'b1110;
	mem[2193] = 4'b1110;
	mem[2194] = 4'b1110;
	mem[2195] = 4'b1110;
	mem[2196] = 4'b1111;
	mem[2197] = 4'b1111;
	mem[2198] = 4'b1111;
	mem[2199] = 4'b1101;
	mem[2200] = 4'b1101;
	mem[2201] = 4'b1101;
	mem[2202] = 4'b1111;
	mem[2203] = 4'b1111;
	mem[2204] = 4'b1111;
	mem[2205] = 4'b1111;
	mem[2206] = 4'b1111;
	mem[2207] = 4'b1101;
	mem[2208] = 4'b1101;
	mem[2209] = 4'b1110;
	mem[2210] = 4'b1111;
	mem[2211] = 4'b1111;
	mem[2212] = 4'b1111;
	mem[2213] = 4'b1001;
	mem[2214] = 4'b0110;
	mem[2215] = 4'b0110;
	mem[2216] = 4'b0110;
	mem[2217] = 4'b0110;
	mem[2218] = 4'b0110;
	mem[2219] = 4'b0110;
	mem[2220] = 4'b0110;
	mem[2221] = 4'b0110;
	mem[2222] = 4'b0110;
	mem[2223] = 4'b0110;
	mem[2224] = 4'b0110;
	mem[2225] = 4'b0110;
	mem[2226] = 4'b0110;
	mem[2227] = 4'b0110;
	mem[2228] = 4'b0111;
	mem[2229] = 4'b0111;
	mem[2230] = 4'b0111;
	mem[2231] = 4'b0111;
	mem[2232] = 4'b0111;
	mem[2233] = 4'b0111;
	mem[2234] = 4'b0111;
	mem[2235] = 4'b0101;
	mem[2236] = 4'b0011;
	mem[2237] = 4'b0001;
	mem[2238] = 4'b0000;
	mem[2239] = 4'b0000;
	mem[2240] = 4'b0000;
	mem[2241] = 4'b0000;
	mem[2242] = 4'b0000;
	mem[2243] = 4'b0000;
	mem[2244] = 4'b0000;
	mem[2245] = 4'b0000;
	mem[2246] = 4'b0000;
	mem[2247] = 4'b1100;
	mem[2248] = 4'b1111;
	mem[2249] = 4'b1111;
	mem[2250] = 4'b1111;
	mem[2251] = 4'b1111;
	mem[2252] = 4'b1111;
	mem[2253] = 4'b1111;
	mem[2254] = 4'b1111;
	mem[2255] = 4'b1111;
	mem[2256] = 4'b1111;
	mem[2257] = 4'b1111;
	mem[2258] = 4'b1111;
	mem[2259] = 4'b1111;
	mem[2260] = 4'b1111;
	mem[2261] = 4'b1111;
	mem[2262] = 4'b1111;
	mem[2263] = 4'b1110;
	mem[2264] = 4'b1101;
	mem[2265] = 4'b1101;
	mem[2266] = 4'b1110;
	mem[2267] = 4'b1111;
	mem[2268] = 4'b1111;
	mem[2269] = 4'b1111;
	mem[2270] = 4'b1111;
	mem[2271] = 4'b1111;
	mem[2272] = 4'b1111;
	mem[2273] = 4'b1111;
	mem[2274] = 4'b1111;
	mem[2275] = 4'b1111;
	mem[2276] = 4'b1111;
	mem[2277] = 4'b1111;
	mem[2278] = 4'b1111;
	mem[2279] = 4'b1111;
	mem[2280] = 4'b1111;
	mem[2281] = 4'b0110;
	mem[2282] = 4'b0000;
	mem[2283] = 4'b0000;
	mem[2284] = 4'b0000;
	mem[2285] = 4'b0000;
	mem[2286] = 4'b0000;
	mem[2287] = 4'b0000;
	mem[2288] = 4'b0000;
	mem[2289] = 4'b0000;
	mem[2290] = 4'b0000;
	mem[2291] = 4'b0000;
	mem[2292] = 4'b0000;
	mem[2293] = 4'b0000;
	mem[2294] = 4'b0000;
	mem[2295] = 4'b0000;
	mem[2296] = 4'b0000;
	mem[2297] = 4'b0000;
	mem[2298] = 4'b0000;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0111;
	mem[2308] = 4'b1100;
	mem[2309] = 4'b1101;
	mem[2310] = 4'b1101;
	mem[2311] = 4'b1101;
	mem[2312] = 4'b1101;
	mem[2313] = 4'b1101;
	mem[2314] = 4'b1101;
	mem[2315] = 4'b1101;
	mem[2316] = 4'b1101;
	mem[2317] = 4'b1101;
	mem[2318] = 4'b1110;
	mem[2319] = 4'b1110;
	mem[2320] = 4'b1110;
	mem[2321] = 4'b1110;
	mem[2322] = 4'b1110;
	mem[2323] = 4'b1110;
	mem[2324] = 4'b1111;
	mem[2325] = 4'b1111;
	mem[2326] = 4'b1111;
	mem[2327] = 4'b1111;
	mem[2328] = 4'b1101;
	mem[2329] = 4'b1101;
	mem[2330] = 4'b1110;
	mem[2331] = 4'b1111;
	mem[2332] = 4'b1111;
	mem[2333] = 4'b1111;
	mem[2334] = 4'b1111;
	mem[2335] = 4'b1111;
	mem[2336] = 4'b1101;
	mem[2337] = 4'b1110;
	mem[2338] = 4'b1111;
	mem[2339] = 4'b1111;
	mem[2340] = 4'b1111;
	mem[2341] = 4'b1001;
	mem[2342] = 4'b0110;
	mem[2343] = 4'b0110;
	mem[2344] = 4'b0110;
	mem[2345] = 4'b0110;
	mem[2346] = 4'b0110;
	mem[2347] = 4'b0110;
	mem[2348] = 4'b0110;
	mem[2349] = 4'b0110;
	mem[2350] = 4'b0110;
	mem[2351] = 4'b0110;
	mem[2352] = 4'b0110;
	mem[2353] = 4'b0110;
	mem[2354] = 4'b0111;
	mem[2355] = 4'b0111;
	mem[2356] = 4'b0111;
	mem[2357] = 4'b0111;
	mem[2358] = 4'b0111;
	mem[2359] = 4'b0111;
	mem[2360] = 4'b0101;
	mem[2361] = 4'b0011;
	mem[2362] = 4'b0001;
	mem[2363] = 4'b0000;
	mem[2364] = 4'b0000;
	mem[2365] = 4'b0000;
	mem[2366] = 4'b0000;
	mem[2367] = 4'b0000;
	mem[2368] = 4'b0000;
	mem[2369] = 4'b0000;
	mem[2370] = 4'b0000;
	mem[2371] = 4'b0000;
	mem[2372] = 4'b0000;
	mem[2373] = 4'b0000;
	mem[2374] = 4'b0000;
	mem[2375] = 4'b1100;
	mem[2376] = 4'b1111;
	mem[2377] = 4'b1111;
	mem[2378] = 4'b1111;
	mem[2379] = 4'b1111;
	mem[2380] = 4'b1111;
	mem[2381] = 4'b1111;
	mem[2382] = 4'b1111;
	mem[2383] = 4'b1111;
	mem[2384] = 4'b1111;
	mem[2385] = 4'b1111;
	mem[2386] = 4'b1111;
	mem[2387] = 4'b1111;
	mem[2388] = 4'b1111;
	mem[2389] = 4'b1111;
	mem[2390] = 4'b1111;
	mem[2391] = 4'b1111;
	mem[2392] = 4'b1111;
	mem[2393] = 4'b1111;
	mem[2394] = 4'b1111;
	mem[2395] = 4'b1111;
	mem[2396] = 4'b1111;
	mem[2397] = 4'b1111;
	mem[2398] = 4'b1111;
	mem[2399] = 4'b1111;
	mem[2400] = 4'b1111;
	mem[2401] = 4'b1111;
	mem[2402] = 4'b1111;
	mem[2403] = 4'b1111;
	mem[2404] = 4'b1111;
	mem[2405] = 4'b1111;
	mem[2406] = 4'b1111;
	mem[2407] = 4'b1111;
	mem[2408] = 4'b1111;
	mem[2409] = 4'b0110;
	mem[2410] = 4'b0000;
	mem[2411] = 4'b0000;
	mem[2412] = 4'b0000;
	mem[2413] = 4'b0000;
	mem[2414] = 4'b0000;
	mem[2415] = 4'b0000;
	mem[2416] = 4'b0000;
	mem[2417] = 4'b0000;
	mem[2418] = 4'b0000;
	mem[2419] = 4'b0000;
	mem[2420] = 4'b0000;
	mem[2421] = 4'b0000;
	mem[2422] = 4'b0000;
	mem[2423] = 4'b0000;
	mem[2424] = 4'b0000;
	mem[2425] = 4'b0000;
	mem[2426] = 4'b0000;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0111;
	mem[2436] = 4'b1100;
	mem[2437] = 4'b1101;
	mem[2438] = 4'b1101;
	mem[2439] = 4'b1101;
	mem[2440] = 4'b1101;
	mem[2441] = 4'b1101;
	mem[2442] = 4'b1101;
	mem[2443] = 4'b1101;
	mem[2444] = 4'b1110;
	mem[2445] = 4'b1110;
	mem[2446] = 4'b1110;
	mem[2447] = 4'b1110;
	mem[2448] = 4'b1110;
	mem[2449] = 4'b1110;
	mem[2450] = 4'b1110;
	mem[2451] = 4'b1110;
	mem[2452] = 4'b1111;
	mem[2453] = 4'b1111;
	mem[2454] = 4'b1111;
	mem[2455] = 4'b1111;
	mem[2456] = 4'b1111;
	mem[2457] = 4'b1101;
	mem[2458] = 4'b1101;
	mem[2459] = 4'b1110;
	mem[2460] = 4'b1111;
	mem[2461] = 4'b1111;
	mem[2462] = 4'b1111;
	mem[2463] = 4'b1111;
	mem[2464] = 4'b1111;
	mem[2465] = 4'b1111;
	mem[2466] = 4'b1111;
	mem[2467] = 4'b1111;
	mem[2468] = 4'b1111;
	mem[2469] = 4'b1001;
	mem[2470] = 4'b0110;
	mem[2471] = 4'b0110;
	mem[2472] = 4'b0110;
	mem[2473] = 4'b0110;
	mem[2474] = 4'b0110;
	mem[2475] = 4'b0110;
	mem[2476] = 4'b0110;
	mem[2477] = 4'b0110;
	mem[2478] = 4'b0110;
	mem[2479] = 4'b0110;
	mem[2480] = 4'b0110;
	mem[2481] = 4'b0111;
	mem[2482] = 4'b0111;
	mem[2483] = 4'b0111;
	mem[2484] = 4'b0111;
	mem[2485] = 4'b0110;
	mem[2486] = 4'b0011;
	mem[2487] = 4'b0001;
	mem[2488] = 4'b0000;
	mem[2489] = 4'b0000;
	mem[2490] = 4'b0000;
	mem[2491] = 4'b0000;
	mem[2492] = 4'b0000;
	mem[2493] = 4'b0000;
	mem[2494] = 4'b0000;
	mem[2495] = 4'b0000;
	mem[2496] = 4'b0000;
	mem[2497] = 4'b0000;
	mem[2498] = 4'b0000;
	mem[2499] = 4'b0000;
	mem[2500] = 4'b0000;
	mem[2501] = 4'b0000;
	mem[2502] = 4'b0000;
	mem[2503] = 4'b1100;
	mem[2504] = 4'b1111;
	mem[2505] = 4'b1111;
	mem[2506] = 4'b1111;
	mem[2507] = 4'b1111;
	mem[2508] = 4'b1111;
	mem[2509] = 4'b1111;
	mem[2510] = 4'b1111;
	mem[2511] = 4'b1111;
	mem[2512] = 4'b1111;
	mem[2513] = 4'b1111;
	mem[2514] = 4'b1111;
	mem[2515] = 4'b1111;
	mem[2516] = 4'b1110;
	mem[2517] = 4'b1111;
	mem[2518] = 4'b1111;
	mem[2519] = 4'b1111;
	mem[2520] = 4'b1111;
	mem[2521] = 4'b1111;
	mem[2522] = 4'b1111;
	mem[2523] = 4'b1111;
	mem[2524] = 4'b1111;
	mem[2525] = 4'b1111;
	mem[2526] = 4'b1111;
	mem[2527] = 4'b1111;
	mem[2528] = 4'b1111;
	mem[2529] = 4'b1111;
	mem[2530] = 4'b1111;
	mem[2531] = 4'b1111;
	mem[2532] = 4'b1111;
	mem[2533] = 4'b1111;
	mem[2534] = 4'b1111;
	mem[2535] = 4'b1111;
	mem[2536] = 4'b1111;
	mem[2537] = 4'b0110;
	mem[2538] = 4'b0000;
	mem[2539] = 4'b0000;
	mem[2540] = 4'b0000;
	mem[2541] = 4'b0000;
	mem[2542] = 4'b0000;
	mem[2543] = 4'b0000;
	mem[2544] = 4'b0000;
	mem[2545] = 4'b0000;
	mem[2546] = 4'b0000;
	mem[2547] = 4'b0000;
	mem[2548] = 4'b0000;
	mem[2549] = 4'b0000;
	mem[2550] = 4'b0000;
	mem[2551] = 4'b0000;
	mem[2552] = 4'b0000;
	mem[2553] = 4'b0000;
	mem[2554] = 4'b0000;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b0111;
	mem[2564] = 4'b1100;
	mem[2565] = 4'b1101;
	mem[2566] = 4'b1101;
	mem[2567] = 4'b1101;
	mem[2568] = 4'b1101;
	mem[2569] = 4'b1101;
	mem[2570] = 4'b1110;
	mem[2571] = 4'b1110;
	mem[2572] = 4'b1110;
	mem[2573] = 4'b1110;
	mem[2574] = 4'b1110;
	mem[2575] = 4'b1110;
	mem[2576] = 4'b1110;
	mem[2577] = 4'b1110;
	mem[2578] = 4'b1101;
	mem[2579] = 4'b1101;
	mem[2580] = 4'b1110;
	mem[2581] = 4'b1110;
	mem[2582] = 4'b1111;
	mem[2583] = 4'b1111;
	mem[2584] = 4'b1111;
	mem[2585] = 4'b1111;
	mem[2586] = 4'b1101;
	mem[2587] = 4'b1101;
	mem[2588] = 4'b1110;
	mem[2589] = 4'b1111;
	mem[2590] = 4'b1111;
	mem[2591] = 4'b1111;
	mem[2592] = 4'b1111;
	mem[2593] = 4'b1111;
	mem[2594] = 4'b1111;
	mem[2595] = 4'b1111;
	mem[2596] = 4'b1111;
	mem[2597] = 4'b1001;
	mem[2598] = 4'b0110;
	mem[2599] = 4'b0110;
	mem[2600] = 4'b0110;
	mem[2601] = 4'b0110;
	mem[2602] = 4'b0110;
	mem[2603] = 4'b0110;
	mem[2604] = 4'b0110;
	mem[2605] = 4'b0110;
	mem[2606] = 4'b0110;
	mem[2607] = 4'b0111;
	mem[2608] = 4'b0111;
	mem[2609] = 4'b0111;
	mem[2610] = 4'b0110;
	mem[2611] = 4'b0100;
	mem[2612] = 4'b0001;
	mem[2613] = 4'b0000;
	mem[2614] = 4'b0000;
	mem[2615] = 4'b0000;
	mem[2616] = 4'b0000;
	mem[2617] = 4'b0000;
	mem[2618] = 4'b0000;
	mem[2619] = 4'b0000;
	mem[2620] = 4'b0000;
	mem[2621] = 4'b0000;
	mem[2622] = 4'b0000;
	mem[2623] = 4'b0000;
	mem[2624] = 4'b0000;
	mem[2625] = 4'b0000;
	mem[2626] = 4'b0000;
	mem[2627] = 4'b0000;
	mem[2628] = 4'b0000;
	mem[2629] = 4'b0000;
	mem[2630] = 4'b0000;
	mem[2631] = 4'b1011;
	mem[2632] = 4'b1111;
	mem[2633] = 4'b1111;
	mem[2634] = 4'b1111;
	mem[2635] = 4'b1111;
	mem[2636] = 4'b1111;
	mem[2637] = 4'b1111;
	mem[2638] = 4'b1111;
	mem[2639] = 4'b1111;
	mem[2640] = 4'b1111;
	mem[2641] = 4'b1111;
	mem[2642] = 4'b1111;
	mem[2643] = 4'b1111;
	mem[2644] = 4'b1101;
	mem[2645] = 4'b1101;
	mem[2646] = 4'b1111;
	mem[2647] = 4'b1111;
	mem[2648] = 4'b1111;
	mem[2649] = 4'b1111;
	mem[2650] = 4'b1111;
	mem[2651] = 4'b1111;
	mem[2652] = 4'b1111;
	mem[2653] = 4'b1111;
	mem[2654] = 4'b1111;
	mem[2655] = 4'b1111;
	mem[2656] = 4'b1111;
	mem[2657] = 4'b1111;
	mem[2658] = 4'b1111;
	mem[2659] = 4'b1111;
	mem[2660] = 4'b1111;
	mem[2661] = 4'b1111;
	mem[2662] = 4'b1111;
	mem[2663] = 4'b1111;
	mem[2664] = 4'b1111;
	mem[2665] = 4'b0110;
	mem[2666] = 4'b0000;
	mem[2667] = 4'b0000;
	mem[2668] = 4'b0000;
	mem[2669] = 4'b0000;
	mem[2670] = 4'b0000;
	mem[2671] = 4'b0000;
	mem[2672] = 4'b0000;
	mem[2673] = 4'b0000;
	mem[2674] = 4'b0000;
	mem[2675] = 4'b0000;
	mem[2676] = 4'b0000;
	mem[2677] = 4'b0000;
	mem[2678] = 4'b0000;
	mem[2679] = 4'b0000;
	mem[2680] = 4'b0000;
	mem[2681] = 4'b0000;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b0111;
	mem[2692] = 4'b1100;
	mem[2693] = 4'b1101;
	mem[2694] = 4'b1101;
	mem[2695] = 4'b1101;
	mem[2696] = 4'b1110;
	mem[2697] = 4'b1110;
	mem[2698] = 4'b1110;
	mem[2699] = 4'b1110;
	mem[2700] = 4'b1110;
	mem[2701] = 4'b1110;
	mem[2702] = 4'b1110;
	mem[2703] = 4'b1110;
	mem[2704] = 4'b1110;
	mem[2705] = 4'b1101;
	mem[2706] = 4'b1100;
	mem[2707] = 4'b1100;
	mem[2708] = 4'b1101;
	mem[2709] = 4'b1101;
	mem[2710] = 4'b1101;
	mem[2711] = 4'b1110;
	mem[2712] = 4'b1111;
	mem[2713] = 4'b1111;
	mem[2714] = 4'b1111;
	mem[2715] = 4'b1101;
	mem[2716] = 4'b1101;
	mem[2717] = 4'b1110;
	mem[2718] = 4'b1111;
	mem[2719] = 4'b1111;
	mem[2720] = 4'b1111;
	mem[2721] = 4'b1111;
	mem[2722] = 4'b1111;
	mem[2723] = 4'b1111;
	mem[2724] = 4'b1111;
	mem[2725] = 4'b1001;
	mem[2726] = 4'b0110;
	mem[2727] = 4'b0110;
	mem[2728] = 4'b0110;
	mem[2729] = 4'b0110;
	mem[2730] = 4'b0110;
	mem[2731] = 4'b0110;
	mem[2732] = 4'b0110;
	mem[2733] = 4'b0111;
	mem[2734] = 4'b0111;
	mem[2735] = 4'b0111;
	mem[2736] = 4'b0101;
	mem[2737] = 4'b0010;
	mem[2738] = 4'b0000;
	mem[2739] = 4'b0000;
	mem[2740] = 4'b0000;
	mem[2741] = 4'b0000;
	mem[2742] = 4'b0000;
	mem[2743] = 4'b0000;
	mem[2744] = 4'b0000;
	mem[2745] = 4'b0000;
	mem[2746] = 4'b0000;
	mem[2747] = 4'b0000;
	mem[2748] = 4'b0000;
	mem[2749] = 4'b0000;
	mem[2750] = 4'b0000;
	mem[2751] = 4'b0000;
	mem[2752] = 4'b0000;
	mem[2753] = 4'b0000;
	mem[2754] = 4'b0000;
	mem[2755] = 4'b0000;
	mem[2756] = 4'b0000;
	mem[2757] = 4'b0000;
	mem[2758] = 4'b0000;
	mem[2759] = 4'b1010;
	mem[2760] = 4'b1111;
	mem[2761] = 4'b1111;
	mem[2762] = 4'b1111;
	mem[2763] = 4'b1111;
	mem[2764] = 4'b1111;
	mem[2765] = 4'b1111;
	mem[2766] = 4'b1111;
	mem[2767] = 4'b1111;
	mem[2768] = 4'b1111;
	mem[2769] = 4'b1111;
	mem[2770] = 4'b1111;
	mem[2771] = 4'b1101;
	mem[2772] = 4'b1101;
	mem[2773] = 4'b1101;
	mem[2774] = 4'b1101;
	mem[2775] = 4'b1111;
	mem[2776] = 4'b1111;
	mem[2777] = 4'b1111;
	mem[2778] = 4'b1111;
	mem[2779] = 4'b1111;
	mem[2780] = 4'b1111;
	mem[2781] = 4'b1111;
	mem[2782] = 4'b1111;
	mem[2783] = 4'b1111;
	mem[2784] = 4'b1111;
	mem[2785] = 4'b1111;
	mem[2786] = 4'b1111;
	mem[2787] = 4'b1111;
	mem[2788] = 4'b1111;
	mem[2789] = 4'b1111;
	mem[2790] = 4'b1111;
	mem[2791] = 4'b1111;
	mem[2792] = 4'b1111;
	mem[2793] = 4'b0110;
	mem[2794] = 4'b0000;
	mem[2795] = 4'b0000;
	mem[2796] = 4'b0000;
	mem[2797] = 4'b0000;
	mem[2798] = 4'b0000;
	mem[2799] = 4'b0000;
	mem[2800] = 4'b0000;
	mem[2801] = 4'b0000;
	mem[2802] = 4'b0000;
	mem[2803] = 4'b0000;
	mem[2804] = 4'b0000;
	mem[2805] = 4'b0000;
	mem[2806] = 4'b0000;
	mem[2807] = 4'b0000;
	mem[2808] = 4'b0000;
	mem[2809] = 4'b0000;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b0111;
	mem[2820] = 4'b1100;
	mem[2821] = 4'b1101;
	mem[2822] = 4'b1101;
	mem[2823] = 4'b1110;
	mem[2824] = 4'b1110;
	mem[2825] = 4'b1110;
	mem[2826] = 4'b1110;
	mem[2827] = 4'b1110;
	mem[2828] = 4'b1110;
	mem[2829] = 4'b1110;
	mem[2830] = 4'b1110;
	mem[2831] = 4'b1110;
	mem[2832] = 4'b1101;
	mem[2833] = 4'b1100;
	mem[2834] = 4'b1100;
	mem[2835] = 4'b1101;
	mem[2836] = 4'b1111;
	mem[2837] = 4'b1111;
	mem[2838] = 4'b1101;
	mem[2839] = 4'b1101;
	mem[2840] = 4'b1110;
	mem[2841] = 4'b1111;
	mem[2842] = 4'b1111;
	mem[2843] = 4'b1111;
	mem[2844] = 4'b1101;
	mem[2845] = 4'b1110;
	mem[2846] = 4'b1111;
	mem[2847] = 4'b1111;
	mem[2848] = 4'b1111;
	mem[2849] = 4'b1111;
	mem[2850] = 4'b1111;
	mem[2851] = 4'b1111;
	mem[2852] = 4'b1111;
	mem[2853] = 4'b1001;
	mem[2854] = 4'b0110;
	mem[2855] = 4'b0110;
	mem[2856] = 4'b0110;
	mem[2857] = 4'b0110;
	mem[2858] = 4'b0110;
	mem[2859] = 4'b0111;
	mem[2860] = 4'b0111;
	mem[2861] = 4'b0110;
	mem[2862] = 4'b0011;
	mem[2863] = 4'b0001;
	mem[2864] = 4'b0000;
	mem[2865] = 4'b0000;
	mem[2866] = 4'b0000;
	mem[2867] = 4'b0000;
	mem[2868] = 4'b0000;
	mem[2869] = 4'b0000;
	mem[2870] = 4'b0000;
	mem[2871] = 4'b0000;
	mem[2872] = 4'b0000;
	mem[2873] = 4'b0000;
	mem[2874] = 4'b0000;
	mem[2875] = 4'b0000;
	mem[2876] = 4'b0000;
	mem[2877] = 4'b0000;
	mem[2878] = 4'b0000;
	mem[2879] = 4'b0000;
	mem[2880] = 4'b0000;
	mem[2881] = 4'b0000;
	mem[2882] = 4'b0000;
	mem[2883] = 4'b0000;
	mem[2884] = 4'b0000;
	mem[2885] = 4'b0000;
	mem[2886] = 4'b0000;
	mem[2887] = 4'b1010;
	mem[2888] = 4'b1101;
	mem[2889] = 4'b1111;
	mem[2890] = 4'b1111;
	mem[2891] = 4'b1111;
	mem[2892] = 4'b1111;
	mem[2893] = 4'b1111;
	mem[2894] = 4'b1111;
	mem[2895] = 4'b1111;
	mem[2896] = 4'b1111;
	mem[2897] = 4'b1111;
	mem[2898] = 4'b1101;
	mem[2899] = 4'b1101;
	mem[2900] = 4'b1101;
	mem[2901] = 4'b1101;
	mem[2902] = 4'b1110;
	mem[2903] = 4'b1111;
	mem[2904] = 4'b1111;
	mem[2905] = 4'b1111;
	mem[2906] = 4'b1111;
	mem[2907] = 4'b1111;
	mem[2908] = 4'b1111;
	mem[2909] = 4'b1111;
	mem[2910] = 4'b1111;
	mem[2911] = 4'b1111;
	mem[2912] = 4'b1111;
	mem[2913] = 4'b1111;
	mem[2914] = 4'b1111;
	mem[2915] = 4'b1111;
	mem[2916] = 4'b1111;
	mem[2917] = 4'b1111;
	mem[2918] = 4'b1111;
	mem[2919] = 4'b1111;
	mem[2920] = 4'b1111;
	mem[2921] = 4'b0110;
	mem[2922] = 4'b0000;
	mem[2923] = 4'b0000;
	mem[2924] = 4'b0000;
	mem[2925] = 4'b0000;
	mem[2926] = 4'b0000;
	mem[2927] = 4'b0000;
	mem[2928] = 4'b0000;
	mem[2929] = 4'b0000;
	mem[2930] = 4'b0000;
	mem[2931] = 4'b0000;
	mem[2932] = 4'b0000;
	mem[2933] = 4'b0000;
	mem[2934] = 4'b0000;
	mem[2935] = 4'b0000;
	mem[2936] = 4'b0000;
	mem[2937] = 4'b0000;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b0111;
	mem[2948] = 4'b1100;
	mem[2949] = 4'b1101;
	mem[2950] = 4'b1110;
	mem[2951] = 4'b1110;
	mem[2952] = 4'b1110;
	mem[2953] = 4'b1110;
	mem[2954] = 4'b1110;
	mem[2955] = 4'b1110;
	mem[2956] = 4'b1110;
	mem[2957] = 4'b1110;
	mem[2958] = 4'b1110;
	mem[2959] = 4'b1110;
	mem[2960] = 4'b1101;
	mem[2961] = 4'b1100;
	mem[2962] = 4'b1100;
	mem[2963] = 4'b1110;
	mem[2964] = 4'b1111;
	mem[2965] = 4'b1111;
	mem[2966] = 4'b1111;
	mem[2967] = 4'b1101;
	mem[2968] = 4'b1101;
	mem[2969] = 4'b1111;
	mem[2970] = 4'b1111;
	mem[2971] = 4'b1111;
	mem[2972] = 4'b1111;
	mem[2973] = 4'b1111;
	mem[2974] = 4'b1111;
	mem[2975] = 4'b1111;
	mem[2976] = 4'b1111;
	mem[2977] = 4'b1111;
	mem[2978] = 4'b1111;
	mem[2979] = 4'b1111;
	mem[2980] = 4'b1111;
	mem[2981] = 4'b1001;
	mem[2982] = 4'b0110;
	mem[2983] = 4'b0110;
	mem[2984] = 4'b0110;
	mem[2985] = 4'b0111;
	mem[2986] = 4'b0111;
	mem[2987] = 4'b0101;
	mem[2988] = 4'b0010;
	mem[2989] = 4'b0000;
	mem[2990] = 4'b0000;
	mem[2991] = 4'b0000;
	mem[2992] = 4'b0000;
	mem[2993] = 4'b0000;
	mem[2994] = 4'b0000;
	mem[2995] = 4'b0000;
	mem[2996] = 4'b0000;
	mem[2997] = 4'b0000;
	mem[2998] = 4'b0000;
	mem[2999] = 4'b0000;
	mem[3000] = 4'b0000;
	mem[3001] = 4'b0000;
	mem[3002] = 4'b0000;
	mem[3003] = 4'b0000;
	mem[3004] = 4'b0000;
	mem[3005] = 4'b0000;
	mem[3006] = 4'b0000;
	mem[3007] = 4'b0000;
	mem[3008] = 4'b0000;
	mem[3009] = 4'b0000;
	mem[3010] = 4'b0000;
	mem[3011] = 4'b0000;
	mem[3012] = 4'b0000;
	mem[3013] = 4'b0000;
	mem[3014] = 4'b0000;
	mem[3015] = 4'b1010;
	mem[3016] = 4'b1101;
	mem[3017] = 4'b1101;
	mem[3018] = 4'b1111;
	mem[3019] = 4'b1111;
	mem[3020] = 4'b1111;
	mem[3021] = 4'b1111;
	mem[3022] = 4'b1111;
	mem[3023] = 4'b1111;
	mem[3024] = 4'b1111;
	mem[3025] = 4'b1101;
	mem[3026] = 4'b1101;
	mem[3027] = 4'b1101;
	mem[3028] = 4'b1101;
	mem[3029] = 4'b1110;
	mem[3030] = 4'b1111;
	mem[3031] = 4'b1111;
	mem[3032] = 4'b1111;
	mem[3033] = 4'b1111;
	mem[3034] = 4'b1111;
	mem[3035] = 4'b1111;
	mem[3036] = 4'b1111;
	mem[3037] = 4'b1111;
	mem[3038] = 4'b1111;
	mem[3039] = 4'b1111;
	mem[3040] = 4'b1111;
	mem[3041] = 4'b1111;
	mem[3042] = 4'b1111;
	mem[3043] = 4'b1111;
	mem[3044] = 4'b1111;
	mem[3045] = 4'b1111;
	mem[3046] = 4'b1111;
	mem[3047] = 4'b1111;
	mem[3048] = 4'b1111;
	mem[3049] = 4'b0110;
	mem[3050] = 4'b0000;
	mem[3051] = 4'b0000;
	mem[3052] = 4'b0000;
	mem[3053] = 4'b0000;
	mem[3054] = 4'b0000;
	mem[3055] = 4'b0000;
	mem[3056] = 4'b0000;
	mem[3057] = 4'b0000;
	mem[3058] = 4'b0000;
	mem[3059] = 4'b0000;
	mem[3060] = 4'b0000;
	mem[3061] = 4'b0000;
	mem[3062] = 4'b0000;
	mem[3063] = 4'b0000;
	mem[3064] = 4'b0000;
	mem[3065] = 4'b0000;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b0111;
	mem[3076] = 4'b1100;
	mem[3077] = 4'b1101;
	mem[3078] = 4'b1110;
	mem[3079] = 4'b1110;
	mem[3080] = 4'b1110;
	mem[3081] = 4'b1110;
	mem[3082] = 4'b1110;
	mem[3083] = 4'b1110;
	mem[3084] = 4'b1110;
	mem[3085] = 4'b1110;
	mem[3086] = 4'b1110;
	mem[3087] = 4'b1110;
	mem[3088] = 4'b1101;
	mem[3089] = 4'b1100;
	mem[3090] = 4'b1101;
	mem[3091] = 4'b1110;
	mem[3092] = 4'b1111;
	mem[3093] = 4'b1111;
	mem[3094] = 4'b1111;
	mem[3095] = 4'b1111;
	mem[3096] = 4'b1101;
	mem[3097] = 4'b1110;
	mem[3098] = 4'b1111;
	mem[3099] = 4'b1111;
	mem[3100] = 4'b1111;
	mem[3101] = 4'b1111;
	mem[3102] = 4'b1111;
	mem[3103] = 4'b1111;
	mem[3104] = 4'b1111;
	mem[3105] = 4'b1111;
	mem[3106] = 4'b1111;
	mem[3107] = 4'b1111;
	mem[3108] = 4'b1111;
	mem[3109] = 4'b1001;
	mem[3110] = 4'b0110;
	mem[3111] = 4'b0111;
	mem[3112] = 4'b0110;
	mem[3113] = 4'b0100;
	mem[3114] = 4'b0001;
	mem[3115] = 4'b0000;
	mem[3116] = 4'b0000;
	mem[3117] = 4'b0000;
	mem[3118] = 4'b0000;
	mem[3119] = 4'b0000;
	mem[3120] = 4'b0000;
	mem[3121] = 4'b0000;
	mem[3122] = 4'b0000;
	mem[3123] = 4'b0000;
	mem[3124] = 4'b0000;
	mem[3125] = 4'b0000;
	mem[3126] = 4'b0000;
	mem[3127] = 4'b0000;
	mem[3128] = 4'b0000;
	mem[3129] = 4'b0000;
	mem[3130] = 4'b0000;
	mem[3131] = 4'b0000;
	mem[3132] = 4'b0000;
	mem[3133] = 4'b0000;
	mem[3134] = 4'b0000;
	mem[3135] = 4'b0000;
	mem[3136] = 4'b0000;
	mem[3137] = 4'b0000;
	mem[3138] = 4'b0000;
	mem[3139] = 4'b0000;
	mem[3140] = 4'b0000;
	mem[3141] = 4'b0000;
	mem[3142] = 4'b0000;
	mem[3143] = 4'b1010;
	mem[3144] = 4'b1101;
	mem[3145] = 4'b1101;
	mem[3146] = 4'b1101;
	mem[3147] = 4'b1111;
	mem[3148] = 4'b1111;
	mem[3149] = 4'b1111;
	mem[3150] = 4'b1111;
	mem[3151] = 4'b1111;
	mem[3152] = 4'b1101;
	mem[3153] = 4'b1101;
	mem[3154] = 4'b1101;
	mem[3155] = 4'b1101;
	mem[3156] = 4'b1110;
	mem[3157] = 4'b1111;
	mem[3158] = 4'b1111;
	mem[3159] = 4'b1111;
	mem[3160] = 4'b1111;
	mem[3161] = 4'b1111;
	mem[3162] = 4'b1111;
	mem[3163] = 4'b1111;
	mem[3164] = 4'b1111;
	mem[3165] = 4'b1111;
	mem[3166] = 4'b1111;
	mem[3167] = 4'b1111;
	mem[3168] = 4'b1111;
	mem[3169] = 4'b1111;
	mem[3170] = 4'b1111;
	mem[3171] = 4'b1111;
	mem[3172] = 4'b1111;
	mem[3173] = 4'b1111;
	mem[3174] = 4'b1111;
	mem[3175] = 4'b1111;
	mem[3176] = 4'b1111;
	mem[3177] = 4'b0110;
	mem[3178] = 4'b0000;
	mem[3179] = 4'b0000;
	mem[3180] = 4'b0000;
	mem[3181] = 4'b0000;
	mem[3182] = 4'b0000;
	mem[3183] = 4'b0000;
	mem[3184] = 4'b0000;
	mem[3185] = 4'b0000;
	mem[3186] = 4'b0000;
	mem[3187] = 4'b0000;
	mem[3188] = 4'b0000;
	mem[3189] = 4'b0000;
	mem[3190] = 4'b0000;
	mem[3191] = 4'b0000;
	mem[3192] = 4'b0000;
	mem[3193] = 4'b0000;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b0111;
	mem[3204] = 4'b1100;
	mem[3205] = 4'b1101;
	mem[3206] = 4'b1110;
	mem[3207] = 4'b1110;
	mem[3208] = 4'b1110;
	mem[3209] = 4'b1110;
	mem[3210] = 4'b1110;
	mem[3211] = 4'b1110;
	mem[3212] = 4'b1110;
	mem[3213] = 4'b1110;
	mem[3214] = 4'b1110;
	mem[3215] = 4'b1110;
	mem[3216] = 4'b1101;
	mem[3217] = 4'b1100;
	mem[3218] = 4'b1100;
	mem[3219] = 4'b1110;
	mem[3220] = 4'b1111;
	mem[3221] = 4'b1111;
	mem[3222] = 4'b1111;
	mem[3223] = 4'b1111;
	mem[3224] = 4'b1101;
	mem[3225] = 4'b1110;
	mem[3226] = 4'b1111;
	mem[3227] = 4'b1111;
	mem[3228] = 4'b1111;
	mem[3229] = 4'b1111;
	mem[3230] = 4'b1111;
	mem[3231] = 4'b1111;
	mem[3232] = 4'b1111;
	mem[3233] = 4'b1111;
	mem[3234] = 4'b1111;
	mem[3235] = 4'b1111;
	mem[3236] = 4'b1111;
	mem[3237] = 4'b1001;
	mem[3238] = 4'b0110;
	mem[3239] = 4'b0100;
	mem[3240] = 4'b0000;
	mem[3241] = 4'b0000;
	mem[3242] = 4'b0000;
	mem[3243] = 4'b0000;
	mem[3244] = 4'b0000;
	mem[3245] = 4'b0000;
	mem[3246] = 4'b0000;
	mem[3247] = 4'b0000;
	mem[3248] = 4'b0000;
	mem[3249] = 4'b0000;
	mem[3250] = 4'b0000;
	mem[3251] = 4'b0000;
	mem[3252] = 4'b0000;
	mem[3253] = 4'b0000;
	mem[3254] = 4'b0000;
	mem[3255] = 4'b0000;
	mem[3256] = 4'b0000;
	mem[3257] = 4'b0000;
	mem[3258] = 4'b0000;
	mem[3259] = 4'b0000;
	mem[3260] = 4'b0000;
	mem[3261] = 4'b0000;
	mem[3262] = 4'b0000;
	mem[3263] = 4'b0000;
	mem[3264] = 4'b0000;
	mem[3265] = 4'b0000;
	mem[3266] = 4'b0000;
	mem[3267] = 4'b0000;
	mem[3268] = 4'b0000;
	mem[3269] = 4'b0000;
	mem[3270] = 4'b0000;
	mem[3271] = 4'b1010;
	mem[3272] = 4'b1101;
	mem[3273] = 4'b1101;
	mem[3274] = 4'b1101;
	mem[3275] = 4'b1101;
	mem[3276] = 4'b1111;
	mem[3277] = 4'b1111;
	mem[3278] = 4'b1111;
	mem[3279] = 4'b1101;
	mem[3280] = 4'b1101;
	mem[3281] = 4'b1101;
	mem[3282] = 4'b1101;
	mem[3283] = 4'b1110;
	mem[3284] = 4'b1111;
	mem[3285] = 4'b1111;
	mem[3286] = 4'b1111;
	mem[3287] = 4'b1111;
	mem[3288] = 4'b1111;
	mem[3289] = 4'b1111;
	mem[3290] = 4'b1111;
	mem[3291] = 4'b1111;
	mem[3292] = 4'b1111;
	mem[3293] = 4'b1111;
	mem[3294] = 4'b1111;
	mem[3295] = 4'b1111;
	mem[3296] = 4'b1111;
	mem[3297] = 4'b1111;
	mem[3298] = 4'b1111;
	mem[3299] = 4'b1111;
	mem[3300] = 4'b1111;
	mem[3301] = 4'b1111;
	mem[3302] = 4'b1111;
	mem[3303] = 4'b1111;
	mem[3304] = 4'b1111;
	mem[3305] = 4'b0110;
	mem[3306] = 4'b0000;
	mem[3307] = 4'b0000;
	mem[3308] = 4'b0000;
	mem[3309] = 4'b0000;
	mem[3310] = 4'b0000;
	mem[3311] = 4'b0000;
	mem[3312] = 4'b0000;
	mem[3313] = 4'b0000;
	mem[3314] = 4'b0000;
	mem[3315] = 4'b0000;
	mem[3316] = 4'b0000;
	mem[3317] = 4'b0000;
	mem[3318] = 4'b0000;
	mem[3319] = 4'b0000;
	mem[3320] = 4'b0000;
	mem[3321] = 4'b0000;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b0111;
	mem[3332] = 4'b1100;
	mem[3333] = 4'b1101;
	mem[3334] = 4'b1110;
	mem[3335] = 4'b1110;
	mem[3336] = 4'b1110;
	mem[3337] = 4'b1110;
	mem[3338] = 4'b1110;
	mem[3339] = 4'b1110;
	mem[3340] = 4'b1110;
	mem[3341] = 4'b1101;
	mem[3342] = 4'b1110;
	mem[3343] = 4'b1110;
	mem[3344] = 4'b1101;
	mem[3345] = 4'b1100;
	mem[3346] = 4'b1100;
	mem[3347] = 4'b1100;
	mem[3348] = 4'b1111;
	mem[3349] = 4'b1111;
	mem[3350] = 4'b1111;
	mem[3351] = 4'b1110;
	mem[3352] = 4'b1101;
	mem[3353] = 4'b1111;
	mem[3354] = 4'b1111;
	mem[3355] = 4'b1111;
	mem[3356] = 4'b1111;
	mem[3357] = 4'b1111;
	mem[3358] = 4'b1111;
	mem[3359] = 4'b1111;
	mem[3360] = 4'b1111;
	mem[3361] = 4'b1111;
	mem[3362] = 4'b1111;
	mem[3363] = 4'b1111;
	mem[3364] = 4'b1111;
	mem[3365] = 4'b0110;
	mem[3366] = 4'b0000;
	mem[3367] = 4'b0000;
	mem[3368] = 4'b0000;
	mem[3369] = 4'b0000;
	mem[3370] = 4'b0000;
	mem[3371] = 4'b0000;
	mem[3372] = 4'b0000;
	mem[3373] = 4'b0000;
	mem[3374] = 4'b0000;
	mem[3375] = 4'b0000;
	mem[3376] = 4'b0000;
	mem[3377] = 4'b0000;
	mem[3378] = 4'b0000;
	mem[3379] = 4'b0000;
	mem[3380] = 4'b0000;
	mem[3381] = 4'b0000;
	mem[3382] = 4'b0000;
	mem[3383] = 4'b0000;
	mem[3384] = 4'b0000;
	mem[3385] = 4'b0000;
	mem[3386] = 4'b0000;
	mem[3387] = 4'b0000;
	mem[3388] = 4'b0000;
	mem[3389] = 4'b0000;
	mem[3390] = 4'b0000;
	mem[3391] = 4'b0000;
	mem[3392] = 4'b0000;
	mem[3393] = 4'b0000;
	mem[3394] = 4'b0000;
	mem[3395] = 4'b0000;
	mem[3396] = 4'b0000;
	mem[3397] = 4'b0000;
	mem[3398] = 4'b0000;
	mem[3399] = 4'b1011;
	mem[3400] = 4'b1101;
	mem[3401] = 4'b1101;
	mem[3402] = 4'b1101;
	mem[3403] = 4'b1101;
	mem[3404] = 4'b1101;
	mem[3405] = 4'b1110;
	mem[3406] = 4'b1101;
	mem[3407] = 4'b1101;
	mem[3408] = 4'b1101;
	mem[3409] = 4'b1101;
	mem[3410] = 4'b1110;
	mem[3411] = 4'b1111;
	mem[3412] = 4'b1111;
	mem[3413] = 4'b1111;
	mem[3414] = 4'b1111;
	mem[3415] = 4'b1111;
	mem[3416] = 4'b1111;
	mem[3417] = 4'b1111;
	mem[3418] = 4'b1111;
	mem[3419] = 4'b1111;
	mem[3420] = 4'b1111;
	mem[3421] = 4'b1111;
	mem[3422] = 4'b1111;
	mem[3423] = 4'b1111;
	mem[3424] = 4'b1111;
	mem[3425] = 4'b1111;
	mem[3426] = 4'b1111;
	mem[3427] = 4'b1111;
	mem[3428] = 4'b1111;
	mem[3429] = 4'b1111;
	mem[3430] = 4'b1111;
	mem[3431] = 4'b1111;
	mem[3432] = 4'b1111;
	mem[3433] = 4'b0110;
	mem[3434] = 4'b0000;
	mem[3435] = 4'b0000;
	mem[3436] = 4'b0000;
	mem[3437] = 4'b0000;
	mem[3438] = 4'b0000;
	mem[3439] = 4'b0000;
	mem[3440] = 4'b0000;
	mem[3441] = 4'b0000;
	mem[3442] = 4'b0000;
	mem[3443] = 4'b0001;
	mem[3444] = 4'b0001;
	mem[3445] = 4'b0000;
	mem[3446] = 4'b0000;
	mem[3447] = 4'b0000;
	mem[3448] = 4'b0000;
	mem[3449] = 4'b0000;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b0111;
	mem[3460] = 4'b1100;
	mem[3461] = 4'b1101;
	mem[3462] = 4'b1110;
	mem[3463] = 4'b1110;
	mem[3464] = 4'b1110;
	mem[3465] = 4'b1110;
	mem[3466] = 4'b1110;
	mem[3467] = 4'b1101;
	mem[3468] = 4'b1100;
	mem[3469] = 4'b1100;
	mem[3470] = 4'b1100;
	mem[3471] = 4'b1101;
	mem[3472] = 4'b1110;
	mem[3473] = 4'b1101;
	mem[3474] = 4'b1100;
	mem[3475] = 4'b1100;
	mem[3476] = 4'b1101;
	mem[3477] = 4'b1110;
	mem[3478] = 4'b1110;
	mem[3479] = 4'b1101;
	mem[3480] = 4'b1110;
	mem[3481] = 4'b1111;
	mem[3482] = 4'b1111;
	mem[3483] = 4'b1111;
	mem[3484] = 4'b1111;
	mem[3485] = 4'b1111;
	mem[3486] = 4'b1111;
	mem[3487] = 4'b1111;
	mem[3488] = 4'b1111;
	mem[3489] = 4'b1111;
	mem[3490] = 4'b1111;
	mem[3491] = 4'b1111;
	mem[3492] = 4'b1111;
	mem[3493] = 4'b0100;
	mem[3494] = 4'b0000;
	mem[3495] = 4'b0000;
	mem[3496] = 4'b0000;
	mem[3497] = 4'b0000;
	mem[3498] = 4'b0000;
	mem[3499] = 4'b0000;
	mem[3500] = 4'b0000;
	mem[3501] = 4'b0000;
	mem[3502] = 4'b0000;
	mem[3503] = 4'b0000;
	mem[3504] = 4'b0000;
	mem[3505] = 4'b0000;
	mem[3506] = 4'b0000;
	mem[3507] = 4'b0000;
	mem[3508] = 4'b0000;
	mem[3509] = 4'b0000;
	mem[3510] = 4'b0000;
	mem[3511] = 4'b0000;
	mem[3512] = 4'b0000;
	mem[3513] = 4'b0000;
	mem[3514] = 4'b0000;
	mem[3515] = 4'b0000;
	mem[3516] = 4'b0000;
	mem[3517] = 4'b0000;
	mem[3518] = 4'b0000;
	mem[3519] = 4'b0000;
	mem[3520] = 4'b0000;
	mem[3521] = 4'b0000;
	mem[3522] = 4'b0000;
	mem[3523] = 4'b0000;
	mem[3524] = 4'b0000;
	mem[3525] = 4'b0000;
	mem[3526] = 4'b0000;
	mem[3527] = 4'b1100;
	mem[3528] = 4'b1111;
	mem[3529] = 4'b1101;
	mem[3530] = 4'b1101;
	mem[3531] = 4'b1101;
	mem[3532] = 4'b1101;
	mem[3533] = 4'b1101;
	mem[3534] = 4'b1101;
	mem[3535] = 4'b1101;
	mem[3536] = 4'b1101;
	mem[3537] = 4'b1110;
	mem[3538] = 4'b1111;
	mem[3539] = 4'b1111;
	mem[3540] = 4'b1111;
	mem[3541] = 4'b1111;
	mem[3542] = 4'b1111;
	mem[3543] = 4'b1111;
	mem[3544] = 4'b1111;
	mem[3545] = 4'b1111;
	mem[3546] = 4'b1111;
	mem[3547] = 4'b1111;
	mem[3548] = 4'b1111;
	mem[3549] = 4'b1111;
	mem[3550] = 4'b1111;
	mem[3551] = 4'b1111;
	mem[3552] = 4'b1111;
	mem[3553] = 4'b1111;
	mem[3554] = 4'b1111;
	mem[3555] = 4'b1111;
	mem[3556] = 4'b1111;
	mem[3557] = 4'b1111;
	mem[3558] = 4'b1111;
	mem[3559] = 4'b1111;
	mem[3560] = 4'b1111;
	mem[3561] = 4'b0110;
	mem[3562] = 4'b0000;
	mem[3563] = 4'b0000;
	mem[3564] = 4'b0000;
	mem[3565] = 4'b0000;
	mem[3566] = 4'b0000;
	mem[3567] = 4'b0000;
	mem[3568] = 4'b0000;
	mem[3569] = 4'b0000;
	mem[3570] = 4'b0001;
	mem[3571] = 4'b0001;
	mem[3572] = 4'b0000;
	mem[3573] = 4'b0000;
	mem[3574] = 4'b0000;
	mem[3575] = 4'b0000;
	mem[3576] = 4'b0000;
	mem[3577] = 4'b0000;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b0111;
	mem[3588] = 4'b1100;
	mem[3589] = 4'b1101;
	mem[3590] = 4'b1110;
	mem[3591] = 4'b1110;
	mem[3592] = 4'b1110;
	mem[3593] = 4'b1110;
	mem[3594] = 4'b1101;
	mem[3595] = 4'b1100;
	mem[3596] = 4'b1100;
	mem[3597] = 4'b1100;
	mem[3598] = 4'b1100;
	mem[3599] = 4'b1110;
	mem[3600] = 4'b1110;
	mem[3601] = 4'b1110;
	mem[3602] = 4'b1101;
	mem[3603] = 4'b1100;
	mem[3604] = 4'b1101;
	mem[3605] = 4'b1101;
	mem[3606] = 4'b1101;
	mem[3607] = 4'b1110;
	mem[3608] = 4'b1111;
	mem[3609] = 4'b1111;
	mem[3610] = 4'b1111;
	mem[3611] = 4'b1111;
	mem[3612] = 4'b1111;
	mem[3613] = 4'b1111;
	mem[3614] = 4'b1111;
	mem[3615] = 4'b1111;
	mem[3616] = 4'b1111;
	mem[3617] = 4'b1111;
	mem[3618] = 4'b1111;
	mem[3619] = 4'b1111;
	mem[3620] = 4'b1111;
	mem[3621] = 4'b0100;
	mem[3622] = 4'b0000;
	mem[3623] = 4'b0000;
	mem[3624] = 4'b0000;
	mem[3625] = 4'b0000;
	mem[3626] = 4'b0000;
	mem[3627] = 4'b0000;
	mem[3628] = 4'b0000;
	mem[3629] = 4'b0000;
	mem[3630] = 4'b0000;
	mem[3631] = 4'b0000;
	mem[3632] = 4'b0000;
	mem[3633] = 4'b0000;
	mem[3634] = 4'b0000;
	mem[3635] = 4'b0000;
	mem[3636] = 4'b0000;
	mem[3637] = 4'b0000;
	mem[3638] = 4'b0000;
	mem[3639] = 4'b0000;
	mem[3640] = 4'b0000;
	mem[3641] = 4'b0000;
	mem[3642] = 4'b0000;
	mem[3643] = 4'b0000;
	mem[3644] = 4'b0000;
	mem[3645] = 4'b0000;
	mem[3646] = 4'b0000;
	mem[3647] = 4'b0000;
	mem[3648] = 4'b0000;
	mem[3649] = 4'b0000;
	mem[3650] = 4'b0000;
	mem[3651] = 4'b0000;
	mem[3652] = 4'b0000;
	mem[3653] = 4'b0000;
	mem[3654] = 4'b0000;
	mem[3655] = 4'b1100;
	mem[3656] = 4'b1111;
	mem[3657] = 4'b1111;
	mem[3658] = 4'b1101;
	mem[3659] = 4'b1101;
	mem[3660] = 4'b1101;
	mem[3661] = 4'b1101;
	mem[3662] = 4'b1101;
	mem[3663] = 4'b1101;
	mem[3664] = 4'b1110;
	mem[3665] = 4'b1111;
	mem[3666] = 4'b1111;
	mem[3667] = 4'b1111;
	mem[3668] = 4'b1111;
	mem[3669] = 4'b1111;
	mem[3670] = 4'b1111;
	mem[3671] = 4'b1111;
	mem[3672] = 4'b1111;
	mem[3673] = 4'b1111;
	mem[3674] = 4'b1111;
	mem[3675] = 4'b1111;
	mem[3676] = 4'b1111;
	mem[3677] = 4'b1111;
	mem[3678] = 4'b1111;
	mem[3679] = 4'b1111;
	mem[3680] = 4'b1111;
	mem[3681] = 4'b1111;
	mem[3682] = 4'b1111;
	mem[3683] = 4'b1111;
	mem[3684] = 4'b1111;
	mem[3685] = 4'b1111;
	mem[3686] = 4'b1111;
	mem[3687] = 4'b1111;
	mem[3688] = 4'b1111;
	mem[3689] = 4'b0110;
	mem[3690] = 4'b0000;
	mem[3691] = 4'b0000;
	mem[3692] = 4'b0000;
	mem[3693] = 4'b0000;
	mem[3694] = 4'b0000;
	mem[3695] = 4'b0000;
	mem[3696] = 4'b0000;
	mem[3697] = 4'b0000;
	mem[3698] = 4'b0001;
	mem[3699] = 4'b0000;
	mem[3700] = 4'b0000;
	mem[3701] = 4'b0000;
	mem[3702] = 4'b0000;
	mem[3703] = 4'b0000;
	mem[3704] = 4'b0000;
	mem[3705] = 4'b0000;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b0111;
	mem[3716] = 4'b1100;
	mem[3717] = 4'b1101;
	mem[3718] = 4'b1110;
	mem[3719] = 4'b1110;
	mem[3720] = 4'b1110;
	mem[3721] = 4'b1101;
	mem[3722] = 4'b1100;
	mem[3723] = 4'b1100;
	mem[3724] = 4'b1101;
	mem[3725] = 4'b1110;
	mem[3726] = 4'b1110;
	mem[3727] = 4'b1110;
	mem[3728] = 4'b1110;
	mem[3729] = 4'b1101;
	mem[3730] = 4'b1110;
	mem[3731] = 4'b1110;
	mem[3732] = 4'b1111;
	mem[3733] = 4'b1111;
	mem[3734] = 4'b1111;
	mem[3735] = 4'b1111;
	mem[3736] = 4'b1111;
	mem[3737] = 4'b1111;
	mem[3738] = 4'b1111;
	mem[3739] = 4'b1111;
	mem[3740] = 4'b1111;
	mem[3741] = 4'b1111;
	mem[3742] = 4'b1111;
	mem[3743] = 4'b1111;
	mem[3744] = 4'b1111;
	mem[3745] = 4'b1111;
	mem[3746] = 4'b1111;
	mem[3747] = 4'b1111;
	mem[3748] = 4'b1111;
	mem[3749] = 4'b0100;
	mem[3750] = 4'b0000;
	mem[3751] = 4'b0000;
	mem[3752] = 4'b0000;
	mem[3753] = 4'b0000;
	mem[3754] = 4'b0000;
	mem[3755] = 4'b0000;
	mem[3756] = 4'b0000;
	mem[3757] = 4'b0000;
	mem[3758] = 4'b0000;
	mem[3759] = 4'b0000;
	mem[3760] = 4'b0000;
	mem[3761] = 4'b0000;
	mem[3762] = 4'b0000;
	mem[3763] = 4'b0000;
	mem[3764] = 4'b0000;
	mem[3765] = 4'b0000;
	mem[3766] = 4'b0000;
	mem[3767] = 4'b0000;
	mem[3768] = 4'b0000;
	mem[3769] = 4'b0000;
	mem[3770] = 4'b0000;
	mem[3771] = 4'b0000;
	mem[3772] = 4'b0000;
	mem[3773] = 4'b0000;
	mem[3774] = 4'b0000;
	mem[3775] = 4'b0000;
	mem[3776] = 4'b0000;
	mem[3777] = 4'b0000;
	mem[3778] = 4'b0000;
	mem[3779] = 4'b0000;
	mem[3780] = 4'b0000;
	mem[3781] = 4'b0000;
	mem[3782] = 4'b0000;
	mem[3783] = 4'b1100;
	mem[3784] = 4'b1111;
	mem[3785] = 4'b1111;
	mem[3786] = 4'b1111;
	mem[3787] = 4'b1101;
	mem[3788] = 4'b1101;
	mem[3789] = 4'b1101;
	mem[3790] = 4'b1101;
	mem[3791] = 4'b1110;
	mem[3792] = 4'b1111;
	mem[3793] = 4'b1111;
	mem[3794] = 4'b1111;
	mem[3795] = 4'b1111;
	mem[3796] = 4'b1111;
	mem[3797] = 4'b1111;
	mem[3798] = 4'b1111;
	mem[3799] = 4'b1111;
	mem[3800] = 4'b1111;
	mem[3801] = 4'b1111;
	mem[3802] = 4'b1111;
	mem[3803] = 4'b1111;
	mem[3804] = 4'b1111;
	mem[3805] = 4'b1111;
	mem[3806] = 4'b1111;
	mem[3807] = 4'b1111;
	mem[3808] = 4'b1111;
	mem[3809] = 4'b1111;
	mem[3810] = 4'b1111;
	mem[3811] = 4'b1111;
	mem[3812] = 4'b1111;
	mem[3813] = 4'b1111;
	mem[3814] = 4'b1111;
	mem[3815] = 4'b1111;
	mem[3816] = 4'b1111;
	mem[3817] = 4'b0110;
	mem[3818] = 4'b0000;
	mem[3819] = 4'b0000;
	mem[3820] = 4'b0000;
	mem[3821] = 4'b0000;
	mem[3822] = 4'b0000;
	mem[3823] = 4'b0000;
	mem[3824] = 4'b0000;
	mem[3825] = 4'b0000;
	mem[3826] = 4'b0000;
	mem[3827] = 4'b0000;
	mem[3828] = 4'b0000;
	mem[3829] = 4'b0000;
	mem[3830] = 4'b0000;
	mem[3831] = 4'b0000;
	mem[3832] = 4'b0000;
	mem[3833] = 4'b0000;
	mem[3834] = 4'b0001;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b0111;
	mem[3844] = 4'b1100;
	mem[3845] = 4'b1101;
	mem[3846] = 4'b1110;
	mem[3847] = 4'b1110;
	mem[3848] = 4'b1110;
	mem[3849] = 4'b1101;
	mem[3850] = 4'b1100;
	mem[3851] = 4'b1100;
	mem[3852] = 4'b1110;
	mem[3853] = 4'b1110;
	mem[3854] = 4'b1110;
	mem[3855] = 4'b1110;
	mem[3856] = 4'b1101;
	mem[3857] = 4'b1100;
	mem[3858] = 4'b1101;
	mem[3859] = 4'b1110;
	mem[3860] = 4'b1111;
	mem[3861] = 4'b1111;
	mem[3862] = 4'b1111;
	mem[3863] = 4'b1111;
	mem[3864] = 4'b1111;
	mem[3865] = 4'b1111;
	mem[3866] = 4'b1111;
	mem[3867] = 4'b1111;
	mem[3868] = 4'b1111;
	mem[3869] = 4'b1111;
	mem[3870] = 4'b1111;
	mem[3871] = 4'b1111;
	mem[3872] = 4'b1111;
	mem[3873] = 4'b1111;
	mem[3874] = 4'b1111;
	mem[3875] = 4'b1111;
	mem[3876] = 4'b1111;
	mem[3877] = 4'b0100;
	mem[3878] = 4'b0000;
	mem[3879] = 4'b0000;
	mem[3880] = 4'b0000;
	mem[3881] = 4'b0000;
	mem[3882] = 4'b0000;
	mem[3883] = 4'b0000;
	mem[3884] = 4'b0000;
	mem[3885] = 4'b0000;
	mem[3886] = 4'b0000;
	mem[3887] = 4'b0000;
	mem[3888] = 4'b0000;
	mem[3889] = 4'b0000;
	mem[3890] = 4'b0000;
	mem[3891] = 4'b0000;
	mem[3892] = 4'b0000;
	mem[3893] = 4'b0000;
	mem[3894] = 4'b0000;
	mem[3895] = 4'b0000;
	mem[3896] = 4'b0000;
	mem[3897] = 4'b0000;
	mem[3898] = 4'b0000;
	mem[3899] = 4'b0000;
	mem[3900] = 4'b0000;
	mem[3901] = 4'b0000;
	mem[3902] = 4'b0000;
	mem[3903] = 4'b0000;
	mem[3904] = 4'b0000;
	mem[3905] = 4'b0000;
	mem[3906] = 4'b0000;
	mem[3907] = 4'b0000;
	mem[3908] = 4'b0000;
	mem[3909] = 4'b0000;
	mem[3910] = 4'b0001;
	mem[3911] = 4'b1100;
	mem[3912] = 4'b1111;
	mem[3913] = 4'b1111;
	mem[3914] = 4'b1111;
	mem[3915] = 4'b1111;
	mem[3916] = 4'b1101;
	mem[3917] = 4'b1101;
	mem[3918] = 4'b1110;
	mem[3919] = 4'b1111;
	mem[3920] = 4'b1111;
	mem[3921] = 4'b1111;
	mem[3922] = 4'b1111;
	mem[3923] = 4'b1111;
	mem[3924] = 4'b1111;
	mem[3925] = 4'b1111;
	mem[3926] = 4'b1111;
	mem[3927] = 4'b1111;
	mem[3928] = 4'b1111;
	mem[3929] = 4'b1111;
	mem[3930] = 4'b1111;
	mem[3931] = 4'b1111;
	mem[3932] = 4'b1111;
	mem[3933] = 4'b1111;
	mem[3934] = 4'b1111;
	mem[3935] = 4'b1111;
	mem[3936] = 4'b1111;
	mem[3937] = 4'b1111;
	mem[3938] = 4'b1111;
	mem[3939] = 4'b1111;
	mem[3940] = 4'b1111;
	mem[3941] = 4'b1111;
	mem[3942] = 4'b1111;
	mem[3943] = 4'b1111;
	mem[3944] = 4'b1111;
	mem[3945] = 4'b0110;
	mem[3946] = 4'b0000;
	mem[3947] = 4'b0000;
	mem[3948] = 4'b0000;
	mem[3949] = 4'b0000;
	mem[3950] = 4'b0000;
	mem[3951] = 4'b0000;
	mem[3952] = 4'b0000;
	mem[3953] = 4'b0000;
	mem[3954] = 4'b0000;
	mem[3955] = 4'b0000;
	mem[3956] = 4'b0000;
	mem[3957] = 4'b0000;
	mem[3958] = 4'b0000;
	mem[3959] = 4'b0000;
	mem[3960] = 4'b0001;
	mem[3961] = 4'b0001;
	mem[3962] = 4'b0001;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b0111;
	mem[3972] = 4'b1011;
	mem[3973] = 4'b1100;
	mem[3974] = 4'b1110;
	mem[3975] = 4'b1110;
	mem[3976] = 4'b1110;
	mem[3977] = 4'b1101;
	mem[3978] = 4'b1100;
	mem[3979] = 4'b1100;
	mem[3980] = 4'b1110;
	mem[3981] = 4'b1110;
	mem[3982] = 4'b1110;
	mem[3983] = 4'b1110;
	mem[3984] = 4'b1101;
	mem[3985] = 4'b1100;
	mem[3986] = 4'b1100;
	mem[3987] = 4'b1110;
	mem[3988] = 4'b1111;
	mem[3989] = 4'b1111;
	mem[3990] = 4'b1111;
	mem[3991] = 4'b1111;
	mem[3992] = 4'b1111;
	mem[3993] = 4'b1111;
	mem[3994] = 4'b1111;
	mem[3995] = 4'b1111;
	mem[3996] = 4'b1111;
	mem[3997] = 4'b1111;
	mem[3998] = 4'b1111;
	mem[3999] = 4'b1111;
	mem[4000] = 4'b1111;
	mem[4001] = 4'b1111;
	mem[4002] = 4'b1111;
	mem[4003] = 4'b1111;
	mem[4004] = 4'b1111;
	mem[4005] = 4'b0100;
	mem[4006] = 4'b0000;
	mem[4007] = 4'b0000;
	mem[4008] = 4'b0000;
	mem[4009] = 4'b0000;
	mem[4010] = 4'b0000;
	mem[4011] = 4'b0000;
	mem[4012] = 4'b0000;
	mem[4013] = 4'b0000;
	mem[4014] = 4'b0000;
	mem[4015] = 4'b0000;
	mem[4016] = 4'b0000;
	mem[4017] = 4'b0000;
	mem[4018] = 4'b0000;
	mem[4019] = 4'b0000;
	mem[4020] = 4'b0000;
	mem[4021] = 4'b0000;
	mem[4022] = 4'b0000;
	mem[4023] = 4'b0000;
	mem[4024] = 4'b0000;
	mem[4025] = 4'b0000;
	mem[4026] = 4'b0000;
	mem[4027] = 4'b0000;
	mem[4028] = 4'b0000;
	mem[4029] = 4'b0000;
	mem[4030] = 4'b0000;
	mem[4031] = 4'b0000;
	mem[4032] = 4'b0000;
	mem[4033] = 4'b0000;
	mem[4034] = 4'b0000;
	mem[4035] = 4'b0000;
	mem[4036] = 4'b0000;
	mem[4037] = 4'b0001;
	mem[4038] = 4'b0000;
	mem[4039] = 4'b1100;
	mem[4040] = 4'b1111;
	mem[4041] = 4'b1111;
	mem[4042] = 4'b1111;
	mem[4043] = 4'b1111;
	mem[4044] = 4'b1111;
	mem[4045] = 4'b1110;
	mem[4046] = 4'b1111;
	mem[4047] = 4'b1111;
	mem[4048] = 4'b1111;
	mem[4049] = 4'b1111;
	mem[4050] = 4'b1111;
	mem[4051] = 4'b1111;
	mem[4052] = 4'b1111;
	mem[4053] = 4'b1111;
	mem[4054] = 4'b1111;
	mem[4055] = 4'b1111;
	mem[4056] = 4'b1111;
	mem[4057] = 4'b1111;
	mem[4058] = 4'b1111;
	mem[4059] = 4'b1111;
	mem[4060] = 4'b1111;
	mem[4061] = 4'b1111;
	mem[4062] = 4'b1111;
	mem[4063] = 4'b1111;
	mem[4064] = 4'b1111;
	mem[4065] = 4'b1111;
	mem[4066] = 4'b1111;
	mem[4067] = 4'b1111;
	mem[4068] = 4'b1111;
	mem[4069] = 4'b1111;
	mem[4070] = 4'b1111;
	mem[4071] = 4'b1111;
	mem[4072] = 4'b1111;
	mem[4073] = 4'b0110;
	mem[4074] = 4'b0000;
	mem[4075] = 4'b0000;
	mem[4076] = 4'b0000;
	mem[4077] = 4'b0000;
	mem[4078] = 4'b0000;
	mem[4079] = 4'b0000;
	mem[4080] = 4'b0000;
	mem[4081] = 4'b0000;
	mem[4082] = 4'b0000;
	mem[4083] = 4'b0000;
	mem[4084] = 4'b0000;
	mem[4085] = 4'b0000;
	mem[4086] = 4'b0000;
	mem[4087] = 4'b0000;
	mem[4088] = 4'b0001;
	mem[4089] = 4'b0000;
	mem[4090] = 4'b0000;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_2r (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0111;
	mem[4] = 4'b1011;
	mem[5] = 4'b1011;
	mem[6] = 4'b1101;
	mem[7] = 4'b1110;
	mem[8] = 4'b1110;
	mem[9] = 4'b1110;
	mem[10] = 4'b1100;
	mem[11] = 4'b1100;
	mem[12] = 4'b1101;
	mem[13] = 4'b1110;
	mem[14] = 4'b1110;
	mem[15] = 4'b1110;
	mem[16] = 4'b1101;
	mem[17] = 4'b1100;
	mem[18] = 4'b1100;
	mem[19] = 4'b1110;
	mem[20] = 4'b1111;
	mem[21] = 4'b1111;
	mem[22] = 4'b1111;
	mem[23] = 4'b1111;
	mem[24] = 4'b1111;
	mem[25] = 4'b1111;
	mem[26] = 4'b1111;
	mem[27] = 4'b1111;
	mem[28] = 4'b1111;
	mem[29] = 4'b1111;
	mem[30] = 4'b1111;
	mem[31] = 4'b1111;
	mem[32] = 4'b1111;
	mem[33] = 4'b1111;
	mem[34] = 4'b1111;
	mem[35] = 4'b1111;
	mem[36] = 4'b1111;
	mem[37] = 4'b0100;
	mem[38] = 4'b0000;
	mem[39] = 4'b0000;
	mem[40] = 4'b0000;
	mem[41] = 4'b0000;
	mem[42] = 4'b0000;
	mem[43] = 4'b0000;
	mem[44] = 4'b0000;
	mem[45] = 4'b0000;
	mem[46] = 4'b0000;
	mem[47] = 4'b0000;
	mem[48] = 4'b0000;
	mem[49] = 4'b0000;
	mem[50] = 4'b0000;
	mem[51] = 4'b0000;
	mem[52] = 4'b0000;
	mem[53] = 4'b0000;
	mem[54] = 4'b0000;
	mem[55] = 4'b0000;
	mem[56] = 4'b0000;
	mem[57] = 4'b0000;
	mem[58] = 4'b0000;
	mem[59] = 4'b0000;
	mem[60] = 4'b0000;
	mem[61] = 4'b0000;
	mem[62] = 4'b0000;
	mem[63] = 4'b0000;
	mem[64] = 4'b0000;
	mem[65] = 4'b0000;
	mem[66] = 4'b0000;
	mem[67] = 4'b0000;
	mem[68] = 4'b0001;
	mem[69] = 4'b0000;
	mem[70] = 4'b0000;
	mem[71] = 4'b1100;
	mem[72] = 4'b1111;
	mem[73] = 4'b1111;
	mem[74] = 4'b1111;
	mem[75] = 4'b1111;
	mem[76] = 4'b1111;
	mem[77] = 4'b1111;
	mem[78] = 4'b1111;
	mem[79] = 4'b1111;
	mem[80] = 4'b1111;
	mem[81] = 4'b1111;
	mem[82] = 4'b1111;
	mem[83] = 4'b1111;
	mem[84] = 4'b1111;
	mem[85] = 4'b1111;
	mem[86] = 4'b1111;
	mem[87] = 4'b1111;
	mem[88] = 4'b1111;
	mem[89] = 4'b1111;
	mem[90] = 4'b1111;
	mem[91] = 4'b1111;
	mem[92] = 4'b1111;
	mem[93] = 4'b1111;
	mem[94] = 4'b1111;
	mem[95] = 4'b1111;
	mem[96] = 4'b1111;
	mem[97] = 4'b1111;
	mem[98] = 4'b1111;
	mem[99] = 4'b1111;
	mem[100] = 4'b1111;
	mem[101] = 4'b1111;
	mem[102] = 4'b1111;
	mem[103] = 4'b1111;
	mem[104] = 4'b1111;
	mem[105] = 4'b0110;
	mem[106] = 4'b0000;
	mem[107] = 4'b0000;
	mem[108] = 4'b0000;
	mem[109] = 4'b0000;
	mem[110] = 4'b0000;
	mem[111] = 4'b0000;
	mem[112] = 4'b0000;
	mem[113] = 4'b0000;
	mem[114] = 4'b0000;
	mem[115] = 4'b0000;
	mem[116] = 4'b0000;
	mem[117] = 4'b0000;
	mem[118] = 4'b0000;
	mem[119] = 4'b0001;
	mem[120] = 4'b0001;
	mem[121] = 4'b0000;
	mem[122] = 4'b0000;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b1000;
	mem[132] = 4'b1100;
	mem[133] = 4'b1011;
	mem[134] = 4'b1100;
	mem[135] = 4'b1101;
	mem[136] = 4'b1110;
	mem[137] = 4'b1110;
	mem[138] = 4'b1101;
	mem[139] = 4'b1100;
	mem[140] = 4'b1100;
	mem[141] = 4'b1101;
	mem[142] = 4'b1101;
	mem[143] = 4'b1101;
	mem[144] = 4'b1100;
	mem[145] = 4'b1100;
	mem[146] = 4'b1101;
	mem[147] = 4'b1110;
	mem[148] = 4'b1111;
	mem[149] = 4'b1111;
	mem[150] = 4'b1111;
	mem[151] = 4'b1111;
	mem[152] = 4'b1111;
	mem[153] = 4'b1111;
	mem[154] = 4'b1111;
	mem[155] = 4'b1111;
	mem[156] = 4'b1111;
	mem[157] = 4'b1111;
	mem[158] = 4'b1111;
	mem[159] = 4'b1111;
	mem[160] = 4'b1111;
	mem[161] = 4'b1111;
	mem[162] = 4'b1111;
	mem[163] = 4'b1111;
	mem[164] = 4'b1111;
	mem[165] = 4'b0100;
	mem[166] = 4'b0000;
	mem[167] = 4'b0000;
	mem[168] = 4'b0000;
	mem[169] = 4'b0000;
	mem[170] = 4'b0000;
	mem[171] = 4'b0000;
	mem[172] = 4'b0000;
	mem[173] = 4'b0000;
	mem[174] = 4'b0000;
	mem[175] = 4'b0000;
	mem[176] = 4'b0000;
	mem[177] = 4'b0000;
	mem[178] = 4'b0000;
	mem[179] = 4'b0000;
	mem[180] = 4'b0000;
	mem[181] = 4'b0000;
	mem[182] = 4'b0000;
	mem[183] = 4'b0000;
	mem[184] = 4'b0000;
	mem[185] = 4'b0000;
	mem[186] = 4'b0000;
	mem[187] = 4'b0000;
	mem[188] = 4'b0000;
	mem[189] = 4'b0000;
	mem[190] = 4'b0000;
	mem[191] = 4'b0000;
	mem[192] = 4'b0000;
	mem[193] = 4'b0000;
	mem[194] = 4'b0000;
	mem[195] = 4'b0001;
	mem[196] = 4'b0000;
	mem[197] = 4'b0000;
	mem[198] = 4'b0000;
	mem[199] = 4'b1100;
	mem[200] = 4'b1111;
	mem[201] = 4'b1111;
	mem[202] = 4'b1111;
	mem[203] = 4'b1111;
	mem[204] = 4'b1111;
	mem[205] = 4'b1111;
	mem[206] = 4'b1111;
	mem[207] = 4'b1111;
	mem[208] = 4'b1111;
	mem[209] = 4'b1111;
	mem[210] = 4'b1111;
	mem[211] = 4'b1111;
	mem[212] = 4'b1111;
	mem[213] = 4'b1111;
	mem[214] = 4'b1111;
	mem[215] = 4'b1111;
	mem[216] = 4'b1111;
	mem[217] = 4'b1111;
	mem[218] = 4'b1111;
	mem[219] = 4'b1111;
	mem[220] = 4'b1111;
	mem[221] = 4'b1111;
	mem[222] = 4'b1111;
	mem[223] = 4'b1111;
	mem[224] = 4'b1111;
	mem[225] = 4'b1111;
	mem[226] = 4'b1111;
	mem[227] = 4'b1111;
	mem[228] = 4'b1111;
	mem[229] = 4'b1111;
	mem[230] = 4'b1111;
	mem[231] = 4'b1111;
	mem[232] = 4'b1111;
	mem[233] = 4'b0110;
	mem[234] = 4'b0000;
	mem[235] = 4'b0000;
	mem[236] = 4'b0000;
	mem[237] = 4'b0000;
	mem[238] = 4'b0000;
	mem[239] = 4'b0000;
	mem[240] = 4'b0000;
	mem[241] = 4'b0000;
	mem[242] = 4'b0000;
	mem[243] = 4'b0000;
	mem[244] = 4'b0001;
	mem[245] = 4'b0001;
	mem[246] = 4'b0001;
	mem[247] = 4'b0001;
	mem[248] = 4'b0000;
	mem[249] = 4'b0000;
	mem[250] = 4'b0000;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0111;
	mem[260] = 4'b1100;
	mem[261] = 4'b1100;
	mem[262] = 4'b1100;
	mem[263] = 4'b1100;
	mem[264] = 4'b1101;
	mem[265] = 4'b1110;
	mem[266] = 4'b1110;
	mem[267] = 4'b1101;
	mem[268] = 4'b1100;
	mem[269] = 4'b1100;
	mem[270] = 4'b1100;
	mem[271] = 4'b1100;
	mem[272] = 4'b1100;
	mem[273] = 4'b1101;
	mem[274] = 4'b1110;
	mem[275] = 4'b1110;
	mem[276] = 4'b1111;
	mem[277] = 4'b1111;
	mem[278] = 4'b1111;
	mem[279] = 4'b1111;
	mem[280] = 4'b1111;
	mem[281] = 4'b1111;
	mem[282] = 4'b1111;
	mem[283] = 4'b1111;
	mem[284] = 4'b1111;
	mem[285] = 4'b1111;
	mem[286] = 4'b1111;
	mem[287] = 4'b1111;
	mem[288] = 4'b1111;
	mem[289] = 4'b1111;
	mem[290] = 4'b1111;
	mem[291] = 4'b1111;
	mem[292] = 4'b1111;
	mem[293] = 4'b0100;
	mem[294] = 4'b0000;
	mem[295] = 4'b0000;
	mem[296] = 4'b0000;
	mem[297] = 4'b0000;
	mem[298] = 4'b0000;
	mem[299] = 4'b0000;
	mem[300] = 4'b0000;
	mem[301] = 4'b0000;
	mem[302] = 4'b0000;
	mem[303] = 4'b0000;
	mem[304] = 4'b0000;
	mem[305] = 4'b0000;
	mem[306] = 4'b0000;
	mem[307] = 4'b0000;
	mem[308] = 4'b0000;
	mem[309] = 4'b0000;
	mem[310] = 4'b0000;
	mem[311] = 4'b0000;
	mem[312] = 4'b0000;
	mem[313] = 4'b0000;
	mem[314] = 4'b0001;
	mem[315] = 4'b0000;
	mem[316] = 4'b0000;
	mem[317] = 4'b0000;
	mem[318] = 4'b0000;
	mem[319] = 4'b0000;
	mem[320] = 4'b0000;
	mem[321] = 4'b0000;
	mem[322] = 4'b0001;
	mem[323] = 4'b0000;
	mem[324] = 4'b0000;
	mem[325] = 4'b0000;
	mem[326] = 4'b0000;
	mem[327] = 4'b1100;
	mem[328] = 4'b1111;
	mem[329] = 4'b1111;
	mem[330] = 4'b1111;
	mem[331] = 4'b1111;
	mem[332] = 4'b1111;
	mem[333] = 4'b1111;
	mem[334] = 4'b1111;
	mem[335] = 4'b1111;
	mem[336] = 4'b1111;
	mem[337] = 4'b1111;
	mem[338] = 4'b1111;
	mem[339] = 4'b1111;
	mem[340] = 4'b1111;
	mem[341] = 4'b1111;
	mem[342] = 4'b1111;
	mem[343] = 4'b1111;
	mem[344] = 4'b1111;
	mem[345] = 4'b1111;
	mem[346] = 4'b1111;
	mem[347] = 4'b1111;
	mem[348] = 4'b1111;
	mem[349] = 4'b1111;
	mem[350] = 4'b1111;
	mem[351] = 4'b1111;
	mem[352] = 4'b1111;
	mem[353] = 4'b1111;
	mem[354] = 4'b1111;
	mem[355] = 4'b1111;
	mem[356] = 4'b1111;
	mem[357] = 4'b1111;
	mem[358] = 4'b1111;
	mem[359] = 4'b1111;
	mem[360] = 4'b1111;
	mem[361] = 4'b0101;
	mem[362] = 4'b0000;
	mem[363] = 4'b0001;
	mem[364] = 4'b0001;
	mem[365] = 4'b0000;
	mem[366] = 4'b0001;
	mem[367] = 4'b0000;
	mem[368] = 4'b0000;
	mem[369] = 4'b0000;
	mem[370] = 4'b0000;
	mem[371] = 4'b0000;
	mem[372] = 4'b0000;
	mem[373] = 4'b0000;
	mem[374] = 4'b0000;
	mem[375] = 4'b0000;
	mem[376] = 4'b0000;
	mem[377] = 4'b0000;
	mem[378] = 4'b0000;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0111;
	mem[388] = 4'b1100;
	mem[389] = 4'b1101;
	mem[390] = 4'b1101;
	mem[391] = 4'b1100;
	mem[392] = 4'b1100;
	mem[393] = 4'b1101;
	mem[394] = 4'b1110;
	mem[395] = 4'b1110;
	mem[396] = 4'b1101;
	mem[397] = 4'b1100;
	mem[398] = 4'b1100;
	mem[399] = 4'b1100;
	mem[400] = 4'b1101;
	mem[401] = 4'b1110;
	mem[402] = 4'b1110;
	mem[403] = 4'b1110;
	mem[404] = 4'b1111;
	mem[405] = 4'b1111;
	mem[406] = 4'b1111;
	mem[407] = 4'b1111;
	mem[408] = 4'b1111;
	mem[409] = 4'b1111;
	mem[410] = 4'b1111;
	mem[411] = 4'b1111;
	mem[412] = 4'b1111;
	mem[413] = 4'b1111;
	mem[414] = 4'b1111;
	mem[415] = 4'b1111;
	mem[416] = 4'b1111;
	mem[417] = 4'b1111;
	mem[418] = 4'b1111;
	mem[419] = 4'b1111;
	mem[420] = 4'b1111;
	mem[421] = 4'b0100;
	mem[422] = 4'b0000;
	mem[423] = 4'b0000;
	mem[424] = 4'b0000;
	mem[425] = 4'b0000;
	mem[426] = 4'b0000;
	mem[427] = 4'b0000;
	mem[428] = 4'b0000;
	mem[429] = 4'b0000;
	mem[430] = 4'b0000;
	mem[431] = 4'b0000;
	mem[432] = 4'b0000;
	mem[433] = 4'b0000;
	mem[434] = 4'b0000;
	mem[435] = 4'b0000;
	mem[436] = 4'b0000;
	mem[437] = 4'b0000;
	mem[438] = 4'b0000;
	mem[439] = 4'b0000;
	mem[440] = 4'b0000;
	mem[441] = 4'b0001;
	mem[442] = 4'b0001;
	mem[443] = 4'b0000;
	mem[444] = 4'b0000;
	mem[445] = 4'b0000;
	mem[446] = 4'b0000;
	mem[447] = 4'b0000;
	mem[448] = 4'b0000;
	mem[449] = 4'b0000;
	mem[450] = 4'b0000;
	mem[451] = 4'b0000;
	mem[452] = 4'b0000;
	mem[453] = 4'b0000;
	mem[454] = 4'b0000;
	mem[455] = 4'b1100;
	mem[456] = 4'b1111;
	mem[457] = 4'b1111;
	mem[458] = 4'b1111;
	mem[459] = 4'b1111;
	mem[460] = 4'b1111;
	mem[461] = 4'b1111;
	mem[462] = 4'b1111;
	mem[463] = 4'b1111;
	mem[464] = 4'b1111;
	mem[465] = 4'b1111;
	mem[466] = 4'b1111;
	mem[467] = 4'b1111;
	mem[468] = 4'b1111;
	mem[469] = 4'b1111;
	mem[470] = 4'b1111;
	mem[471] = 4'b1111;
	mem[472] = 4'b1111;
	mem[473] = 4'b1111;
	mem[474] = 4'b1111;
	mem[475] = 4'b1111;
	mem[476] = 4'b1111;
	mem[477] = 4'b1111;
	mem[478] = 4'b1111;
	mem[479] = 4'b1111;
	mem[480] = 4'b1111;
	mem[481] = 4'b1111;
	mem[482] = 4'b1111;
	mem[483] = 4'b1111;
	mem[484] = 4'b1111;
	mem[485] = 4'b1111;
	mem[486] = 4'b1111;
	mem[487] = 4'b1111;
	mem[488] = 4'b1110;
	mem[489] = 4'b0101;
	mem[490] = 4'b0000;
	mem[491] = 4'b0001;
	mem[492] = 4'b0000;
	mem[493] = 4'b0000;
	mem[494] = 4'b0000;
	mem[495] = 4'b0000;
	mem[496] = 4'b0000;
	mem[497] = 4'b0000;
	mem[498] = 4'b0000;
	mem[499] = 4'b0000;
	mem[500] = 4'b0000;
	mem[501] = 4'b0000;
	mem[502] = 4'b0000;
	mem[503] = 4'b0000;
	mem[504] = 4'b0000;
	mem[505] = 4'b0000;
	mem[506] = 4'b0000;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0111;
	mem[516] = 4'b1100;
	mem[517] = 4'b1101;
	mem[518] = 4'b1110;
	mem[519] = 4'b1101;
	mem[520] = 4'b1100;
	mem[521] = 4'b1100;
	mem[522] = 4'b1101;
	mem[523] = 4'b1110;
	mem[524] = 4'b1110;
	mem[525] = 4'b1110;
	mem[526] = 4'b1110;
	mem[527] = 4'b1110;
	mem[528] = 4'b1110;
	mem[529] = 4'b1110;
	mem[530] = 4'b1110;
	mem[531] = 4'b1101;
	mem[532] = 4'b1111;
	mem[533] = 4'b1111;
	mem[534] = 4'b1111;
	mem[535] = 4'b1111;
	mem[536] = 4'b1111;
	mem[537] = 4'b1111;
	mem[538] = 4'b1111;
	mem[539] = 4'b1111;
	mem[540] = 4'b1111;
	mem[541] = 4'b1111;
	mem[542] = 4'b1111;
	mem[543] = 4'b1111;
	mem[544] = 4'b1111;
	mem[545] = 4'b1111;
	mem[546] = 4'b1111;
	mem[547] = 4'b1111;
	mem[548] = 4'b1111;
	mem[549] = 4'b0100;
	mem[550] = 4'b0000;
	mem[551] = 4'b0000;
	mem[552] = 4'b0000;
	mem[553] = 4'b0000;
	mem[554] = 4'b0000;
	mem[555] = 4'b0000;
	mem[556] = 4'b0000;
	mem[557] = 4'b0000;
	mem[558] = 4'b0000;
	mem[559] = 4'b0000;
	mem[560] = 4'b0000;
	mem[561] = 4'b0000;
	mem[562] = 4'b0000;
	mem[563] = 4'b0000;
	mem[564] = 4'b0000;
	mem[565] = 4'b0000;
	mem[566] = 4'b0001;
	mem[567] = 4'b0001;
	mem[568] = 4'b0001;
	mem[569] = 4'b0001;
	mem[570] = 4'b0000;
	mem[571] = 4'b0000;
	mem[572] = 4'b0000;
	mem[573] = 4'b0000;
	mem[574] = 4'b0000;
	mem[575] = 4'b0000;
	mem[576] = 4'b0000;
	mem[577] = 4'b0000;
	mem[578] = 4'b0000;
	mem[579] = 4'b0000;
	mem[580] = 4'b0000;
	mem[581] = 4'b0000;
	mem[582] = 4'b0000;
	mem[583] = 4'b1100;
	mem[584] = 4'b1111;
	mem[585] = 4'b1111;
	mem[586] = 4'b1111;
	mem[587] = 4'b1111;
	mem[588] = 4'b1111;
	mem[589] = 4'b1111;
	mem[590] = 4'b1111;
	mem[591] = 4'b1111;
	mem[592] = 4'b1111;
	mem[593] = 4'b1111;
	mem[594] = 4'b1111;
	mem[595] = 4'b1111;
	mem[596] = 4'b1111;
	mem[597] = 4'b1111;
	mem[598] = 4'b1111;
	mem[599] = 4'b1111;
	mem[600] = 4'b1111;
	mem[601] = 4'b1111;
	mem[602] = 4'b1111;
	mem[603] = 4'b1111;
	mem[604] = 4'b1111;
	mem[605] = 4'b1111;
	mem[606] = 4'b1111;
	mem[607] = 4'b1111;
	mem[608] = 4'b1111;
	mem[609] = 4'b1111;
	mem[610] = 4'b1111;
	mem[611] = 4'b1111;
	mem[612] = 4'b1111;
	mem[613] = 4'b1111;
	mem[614] = 4'b1111;
	mem[615] = 4'b1111;
	mem[616] = 4'b1111;
	mem[617] = 4'b0101;
	mem[618] = 4'b0000;
	mem[619] = 4'b0000;
	mem[620] = 4'b0000;
	mem[621] = 4'b0000;
	mem[622] = 4'b0000;
	mem[623] = 4'b0000;
	mem[624] = 4'b0000;
	mem[625] = 4'b0000;
	mem[626] = 4'b0000;
	mem[627] = 4'b0001;
	mem[628] = 4'b0000;
	mem[629] = 4'b0000;
	mem[630] = 4'b0000;
	mem[631] = 4'b0000;
	mem[632] = 4'b0000;
	mem[633] = 4'b0000;
	mem[634] = 4'b0000;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0111;
	mem[644] = 4'b1100;
	mem[645] = 4'b1101;
	mem[646] = 4'b1110;
	mem[647] = 4'b1110;
	mem[648] = 4'b1101;
	mem[649] = 4'b1100;
	mem[650] = 4'b1100;
	mem[651] = 4'b1101;
	mem[652] = 4'b1110;
	mem[653] = 4'b1110;
	mem[654] = 4'b1110;
	mem[655] = 4'b1110;
	mem[656] = 4'b1110;
	mem[657] = 4'b1101;
	mem[658] = 4'b1100;
	mem[659] = 4'b1100;
	mem[660] = 4'b1111;
	mem[661] = 4'b1111;
	mem[662] = 4'b1111;
	mem[663] = 4'b1111;
	mem[664] = 4'b1111;
	mem[665] = 4'b1111;
	mem[666] = 4'b1111;
	mem[667] = 4'b1111;
	mem[668] = 4'b1111;
	mem[669] = 4'b1111;
	mem[670] = 4'b1111;
	mem[671] = 4'b1111;
	mem[672] = 4'b1111;
	mem[673] = 4'b1111;
	mem[674] = 4'b1111;
	mem[675] = 4'b1111;
	mem[676] = 4'b1111;
	mem[677] = 4'b0100;
	mem[678] = 4'b0000;
	mem[679] = 4'b0000;
	mem[680] = 4'b0000;
	mem[681] = 4'b0000;
	mem[682] = 4'b0000;
	mem[683] = 4'b0000;
	mem[684] = 4'b0000;
	mem[685] = 4'b0000;
	mem[686] = 4'b0000;
	mem[687] = 4'b0000;
	mem[688] = 4'b0000;
	mem[689] = 4'b0000;
	mem[690] = 4'b0000;
	mem[691] = 4'b0000;
	mem[692] = 4'b0000;
	mem[693] = 4'b0001;
	mem[694] = 4'b0001;
	mem[695] = 4'b0000;
	mem[696] = 4'b0000;
	mem[697] = 4'b0000;
	mem[698] = 4'b0000;
	mem[699] = 4'b0000;
	mem[700] = 4'b0000;
	mem[701] = 4'b0000;
	mem[702] = 4'b0000;
	mem[703] = 4'b0000;
	mem[704] = 4'b0000;
	mem[705] = 4'b0000;
	mem[706] = 4'b0000;
	mem[707] = 4'b0000;
	mem[708] = 4'b0000;
	mem[709] = 4'b0000;
	mem[710] = 4'b0000;
	mem[711] = 4'b1100;
	mem[712] = 4'b1111;
	mem[713] = 4'b1111;
	mem[714] = 4'b1111;
	mem[715] = 4'b1111;
	mem[716] = 4'b1111;
	mem[717] = 4'b1111;
	mem[718] = 4'b1111;
	mem[719] = 4'b1111;
	mem[720] = 4'b1111;
	mem[721] = 4'b1111;
	mem[722] = 4'b1111;
	mem[723] = 4'b1111;
	mem[724] = 4'b1111;
	mem[725] = 4'b1111;
	mem[726] = 4'b1111;
	mem[727] = 4'b1111;
	mem[728] = 4'b1111;
	mem[729] = 4'b1111;
	mem[730] = 4'b1111;
	mem[731] = 4'b1111;
	mem[732] = 4'b1111;
	mem[733] = 4'b1111;
	mem[734] = 4'b1111;
	mem[735] = 4'b1111;
	mem[736] = 4'b1111;
	mem[737] = 4'b1111;
	mem[738] = 4'b1111;
	mem[739] = 4'b1111;
	mem[740] = 4'b1111;
	mem[741] = 4'b1111;
	mem[742] = 4'b1111;
	mem[743] = 4'b1111;
	mem[744] = 4'b1111;
	mem[745] = 4'b0110;
	mem[746] = 4'b0000;
	mem[747] = 4'b0000;
	mem[748] = 4'b0000;
	mem[749] = 4'b0000;
	mem[750] = 4'b0000;
	mem[751] = 4'b0000;
	mem[752] = 4'b0000;
	mem[753] = 4'b0000;
	mem[754] = 4'b0001;
	mem[755] = 4'b0001;
	mem[756] = 4'b0000;
	mem[757] = 4'b0000;
	mem[758] = 4'b0000;
	mem[759] = 4'b0000;
	mem[760] = 4'b0000;
	mem[761] = 4'b0000;
	mem[762] = 4'b0000;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0111;
	mem[772] = 4'b1100;
	mem[773] = 4'b1101;
	mem[774] = 4'b1110;
	mem[775] = 4'b1110;
	mem[776] = 4'b1110;
	mem[777] = 4'b1101;
	mem[778] = 4'b1100;
	mem[779] = 4'b1100;
	mem[780] = 4'b1101;
	mem[781] = 4'b1110;
	mem[782] = 4'b1110;
	mem[783] = 4'b1110;
	mem[784] = 4'b1101;
	mem[785] = 4'b1100;
	mem[786] = 4'b1100;
	mem[787] = 4'b1100;
	mem[788] = 4'b1111;
	mem[789] = 4'b1111;
	mem[790] = 4'b1111;
	mem[791] = 4'b1111;
	mem[792] = 4'b1111;
	mem[793] = 4'b1111;
	mem[794] = 4'b1111;
	mem[795] = 4'b1111;
	mem[796] = 4'b1111;
	mem[797] = 4'b1111;
	mem[798] = 4'b1111;
	mem[799] = 4'b1111;
	mem[800] = 4'b1111;
	mem[801] = 4'b1111;
	mem[802] = 4'b1111;
	mem[803] = 4'b1111;
	mem[804] = 4'b1111;
	mem[805] = 4'b0100;
	mem[806] = 4'b0000;
	mem[807] = 4'b0000;
	mem[808] = 4'b0000;
	mem[809] = 4'b0000;
	mem[810] = 4'b0000;
	mem[811] = 4'b0000;
	mem[812] = 4'b0000;
	mem[813] = 4'b0000;
	mem[814] = 4'b0000;
	mem[815] = 4'b0000;
	mem[816] = 4'b0000;
	mem[817] = 4'b0000;
	mem[818] = 4'b0000;
	mem[819] = 4'b0000;
	mem[820] = 4'b0001;
	mem[821] = 4'b0001;
	mem[822] = 4'b0000;
	mem[823] = 4'b0000;
	mem[824] = 4'b0000;
	mem[825] = 4'b0000;
	mem[826] = 4'b0000;
	mem[827] = 4'b0000;
	mem[828] = 4'b0000;
	mem[829] = 4'b0000;
	mem[830] = 4'b0000;
	mem[831] = 4'b0000;
	mem[832] = 4'b0000;
	mem[833] = 4'b0000;
	mem[834] = 4'b0000;
	mem[835] = 4'b0000;
	mem[836] = 4'b0000;
	mem[837] = 4'b0000;
	mem[838] = 4'b0000;
	mem[839] = 4'b1100;
	mem[840] = 4'b1111;
	mem[841] = 4'b1111;
	mem[842] = 4'b1111;
	mem[843] = 4'b1111;
	mem[844] = 4'b1111;
	mem[845] = 4'b1111;
	mem[846] = 4'b1111;
	mem[847] = 4'b1111;
	mem[848] = 4'b1111;
	mem[849] = 4'b1111;
	mem[850] = 4'b1111;
	mem[851] = 4'b1111;
	mem[852] = 4'b1111;
	mem[853] = 4'b1111;
	mem[854] = 4'b1111;
	mem[855] = 4'b1111;
	mem[856] = 4'b1111;
	mem[857] = 4'b1111;
	mem[858] = 4'b1111;
	mem[859] = 4'b1111;
	mem[860] = 4'b1111;
	mem[861] = 4'b1111;
	mem[862] = 4'b1111;
	mem[863] = 4'b1111;
	mem[864] = 4'b1111;
	mem[865] = 4'b1111;
	mem[866] = 4'b1111;
	mem[867] = 4'b1111;
	mem[868] = 4'b1111;
	mem[869] = 4'b1111;
	mem[870] = 4'b1110;
	mem[871] = 4'b1111;
	mem[872] = 4'b1111;
	mem[873] = 4'b0110;
	mem[874] = 4'b0000;
	mem[875] = 4'b0000;
	mem[876] = 4'b0000;
	mem[877] = 4'b0000;
	mem[878] = 4'b0000;
	mem[879] = 4'b0000;
	mem[880] = 4'b0000;
	mem[881] = 4'b0000;
	mem[882] = 4'b0000;
	mem[883] = 4'b0000;
	mem[884] = 4'b0000;
	mem[885] = 4'b0000;
	mem[886] = 4'b0000;
	mem[887] = 4'b0000;
	mem[888] = 4'b0000;
	mem[889] = 4'b0000;
	mem[890] = 4'b0000;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0111;
	mem[900] = 4'b1100;
	mem[901] = 4'b1101;
	mem[902] = 4'b1110;
	mem[903] = 4'b1110;
	mem[904] = 4'b1110;
	mem[905] = 4'b1110;
	mem[906] = 4'b1101;
	mem[907] = 4'b1100;
	mem[908] = 4'b1101;
	mem[909] = 4'b1110;
	mem[910] = 4'b1101;
	mem[911] = 4'b1101;
	mem[912] = 4'b1100;
	mem[913] = 4'b1100;
	mem[914] = 4'b1100;
	mem[915] = 4'b1100;
	mem[916] = 4'b1111;
	mem[917] = 4'b1111;
	mem[918] = 4'b1111;
	mem[919] = 4'b1111;
	mem[920] = 4'b1111;
	mem[921] = 4'b1111;
	mem[922] = 4'b1111;
	mem[923] = 4'b1111;
	mem[924] = 4'b1111;
	mem[925] = 4'b1111;
	mem[926] = 4'b1111;
	mem[927] = 4'b1111;
	mem[928] = 4'b1111;
	mem[929] = 4'b1111;
	mem[930] = 4'b1111;
	mem[931] = 4'b1111;
	mem[932] = 4'b1111;
	mem[933] = 4'b0100;
	mem[934] = 4'b0000;
	mem[935] = 4'b0000;
	mem[936] = 4'b0000;
	mem[937] = 4'b0000;
	mem[938] = 4'b0000;
	mem[939] = 4'b0000;
	mem[940] = 4'b0000;
	mem[941] = 4'b0000;
	mem[942] = 4'b0000;
	mem[943] = 4'b0000;
	mem[944] = 4'b0000;
	mem[945] = 4'b0000;
	mem[946] = 4'b0000;
	mem[947] = 4'b0000;
	mem[948] = 4'b0001;
	mem[949] = 4'b0000;
	mem[950] = 4'b0000;
	mem[951] = 4'b0000;
	mem[952] = 4'b0000;
	mem[953] = 4'b0000;
	mem[954] = 4'b0000;
	mem[955] = 4'b0000;
	mem[956] = 4'b0000;
	mem[957] = 4'b0000;
	mem[958] = 4'b0000;
	mem[959] = 4'b0000;
	mem[960] = 4'b0000;
	mem[961] = 4'b0001;
	mem[962] = 4'b0000;
	mem[963] = 4'b0000;
	mem[964] = 4'b0000;
	mem[965] = 4'b0000;
	mem[966] = 4'b0000;
	mem[967] = 4'b1100;
	mem[968] = 4'b1111;
	mem[969] = 4'b1111;
	mem[970] = 4'b1111;
	mem[971] = 4'b1111;
	mem[972] = 4'b1111;
	mem[973] = 4'b1111;
	mem[974] = 4'b1111;
	mem[975] = 4'b1111;
	mem[976] = 4'b1111;
	mem[977] = 4'b1111;
	mem[978] = 4'b1111;
	mem[979] = 4'b1111;
	mem[980] = 4'b1111;
	mem[981] = 4'b1111;
	mem[982] = 4'b1111;
	mem[983] = 4'b1111;
	mem[984] = 4'b1111;
	mem[985] = 4'b1111;
	mem[986] = 4'b1111;
	mem[987] = 4'b1111;
	mem[988] = 4'b1111;
	mem[989] = 4'b1111;
	mem[990] = 4'b1111;
	mem[991] = 4'b1111;
	mem[992] = 4'b1111;
	mem[993] = 4'b1111;
	mem[994] = 4'b1111;
	mem[995] = 4'b1111;
	mem[996] = 4'b1110;
	mem[997] = 4'b1101;
	mem[998] = 4'b1101;
	mem[999] = 4'b1101;
	mem[1000] = 4'b1111;
	mem[1001] = 4'b0110;
	mem[1002] = 4'b0000;
	mem[1003] = 4'b0000;
	mem[1004] = 4'b0000;
	mem[1005] = 4'b0000;
	mem[1006] = 4'b0000;
	mem[1007] = 4'b0000;
	mem[1008] = 4'b0000;
	mem[1009] = 4'b0000;
	mem[1010] = 4'b0000;
	mem[1011] = 4'b0000;
	mem[1012] = 4'b0000;
	mem[1013] = 4'b0000;
	mem[1014] = 4'b0000;
	mem[1015] = 4'b0000;
	mem[1016] = 4'b0000;
	mem[1017] = 4'b0000;
	mem[1018] = 4'b0000;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0111;
	mem[1028] = 4'b1100;
	mem[1029] = 4'b1101;
	mem[1030] = 4'b1110;
	mem[1031] = 4'b1110;
	mem[1032] = 4'b1110;
	mem[1033] = 4'b1110;
	mem[1034] = 4'b1110;
	mem[1035] = 4'b1101;
	mem[1036] = 4'b1110;
	mem[1037] = 4'b1101;
	mem[1038] = 4'b1100;
	mem[1039] = 4'b1100;
	mem[1040] = 4'b1100;
	mem[1041] = 4'b1100;
	mem[1042] = 4'b1100;
	mem[1043] = 4'b1100;
	mem[1044] = 4'b1111;
	mem[1045] = 4'b1111;
	mem[1046] = 4'b1111;
	mem[1047] = 4'b1111;
	mem[1048] = 4'b1111;
	mem[1049] = 4'b1111;
	mem[1050] = 4'b1111;
	mem[1051] = 4'b1111;
	mem[1052] = 4'b1111;
	mem[1053] = 4'b1111;
	mem[1054] = 4'b1111;
	mem[1055] = 4'b1111;
	mem[1056] = 4'b1111;
	mem[1057] = 4'b1111;
	mem[1058] = 4'b1111;
	mem[1059] = 4'b1111;
	mem[1060] = 4'b1111;
	mem[1061] = 4'b0100;
	mem[1062] = 4'b0000;
	mem[1063] = 4'b0000;
	mem[1064] = 4'b0000;
	mem[1065] = 4'b0000;
	mem[1066] = 4'b0000;
	mem[1067] = 4'b0000;
	mem[1068] = 4'b0000;
	mem[1069] = 4'b0000;
	mem[1070] = 4'b0000;
	mem[1071] = 4'b0000;
	mem[1072] = 4'b0000;
	mem[1073] = 4'b0000;
	mem[1074] = 4'b0000;
	mem[1075] = 4'b0000;
	mem[1076] = 4'b0000;
	mem[1077] = 4'b0000;
	mem[1078] = 4'b0000;
	mem[1079] = 4'b0000;
	mem[1080] = 4'b0000;
	mem[1081] = 4'b0000;
	mem[1082] = 4'b0000;
	mem[1083] = 4'b0000;
	mem[1084] = 4'b0001;
	mem[1085] = 4'b0000;
	mem[1086] = 4'b0000;
	mem[1087] = 4'b0000;
	mem[1088] = 4'b0000;
	mem[1089] = 4'b0001;
	mem[1090] = 4'b0000;
	mem[1091] = 4'b0000;
	mem[1092] = 4'b0000;
	mem[1093] = 4'b0000;
	mem[1094] = 4'b0000;
	mem[1095] = 4'b1100;
	mem[1096] = 4'b1111;
	mem[1097] = 4'b1111;
	mem[1098] = 4'b1111;
	mem[1099] = 4'b1111;
	mem[1100] = 4'b1111;
	mem[1101] = 4'b1111;
	mem[1102] = 4'b1111;
	mem[1103] = 4'b1111;
	mem[1104] = 4'b1111;
	mem[1105] = 4'b1111;
	mem[1106] = 4'b1111;
	mem[1107] = 4'b1111;
	mem[1108] = 4'b1111;
	mem[1109] = 4'b1111;
	mem[1110] = 4'b1111;
	mem[1111] = 4'b1111;
	mem[1112] = 4'b1111;
	mem[1113] = 4'b1111;
	mem[1114] = 4'b1111;
	mem[1115] = 4'b1111;
	mem[1116] = 4'b1111;
	mem[1117] = 4'b1111;
	mem[1118] = 4'b1111;
	mem[1119] = 4'b1111;
	mem[1120] = 4'b1111;
	mem[1121] = 4'b1111;
	mem[1122] = 4'b1111;
	mem[1123] = 4'b1110;
	mem[1124] = 4'b1101;
	mem[1125] = 4'b1110;
	mem[1126] = 4'b1110;
	mem[1127] = 4'b1101;
	mem[1128] = 4'b1101;
	mem[1129] = 4'b0110;
	mem[1130] = 4'b0000;
	mem[1131] = 4'b0000;
	mem[1132] = 4'b0000;
	mem[1133] = 4'b0000;
	mem[1134] = 4'b0000;
	mem[1135] = 4'b0001;
	mem[1136] = 4'b0000;
	mem[1137] = 4'b0000;
	mem[1138] = 4'b0000;
	mem[1139] = 4'b0000;
	mem[1140] = 4'b0000;
	mem[1141] = 4'b0000;
	mem[1142] = 4'b0000;
	mem[1143] = 4'b0000;
	mem[1144] = 4'b0000;
	mem[1145] = 4'b0000;
	mem[1146] = 4'b0000;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0111;
	mem[1156] = 4'b1100;
	mem[1157] = 4'b1101;
	mem[1158] = 4'b1110;
	mem[1159] = 4'b1110;
	mem[1160] = 4'b1110;
	mem[1161] = 4'b1110;
	mem[1162] = 4'b1110;
	mem[1163] = 4'b1110;
	mem[1164] = 4'b1101;
	mem[1165] = 4'b1100;
	mem[1166] = 4'b1100;
	mem[1167] = 4'b1100;
	mem[1168] = 4'b1100;
	mem[1169] = 4'b1100;
	mem[1170] = 4'b1100;
	mem[1171] = 4'b1100;
	mem[1172] = 4'b1111;
	mem[1173] = 4'b1111;
	mem[1174] = 4'b1111;
	mem[1175] = 4'b1111;
	mem[1176] = 4'b1111;
	mem[1177] = 4'b1111;
	mem[1178] = 4'b1111;
	mem[1179] = 4'b1111;
	mem[1180] = 4'b1111;
	mem[1181] = 4'b1111;
	mem[1182] = 4'b1111;
	mem[1183] = 4'b1111;
	mem[1184] = 4'b1111;
	mem[1185] = 4'b1111;
	mem[1186] = 4'b1111;
	mem[1187] = 4'b1111;
	mem[1188] = 4'b1111;
	mem[1189] = 4'b0100;
	mem[1190] = 4'b0000;
	mem[1191] = 4'b0000;
	mem[1192] = 4'b0000;
	mem[1193] = 4'b0000;
	mem[1194] = 4'b0000;
	mem[1195] = 4'b0000;
	mem[1196] = 4'b0000;
	mem[1197] = 4'b0000;
	mem[1198] = 4'b0000;
	mem[1199] = 4'b0000;
	mem[1200] = 4'b0000;
	mem[1201] = 4'b0000;
	mem[1202] = 4'b0000;
	mem[1203] = 4'b0000;
	mem[1204] = 4'b0000;
	mem[1205] = 4'b0000;
	mem[1206] = 4'b0000;
	mem[1207] = 4'b0000;
	mem[1208] = 4'b0000;
	mem[1209] = 4'b0000;
	mem[1210] = 4'b0000;
	mem[1211] = 4'b0001;
	mem[1212] = 4'b0001;
	mem[1213] = 4'b0000;
	mem[1214] = 4'b0000;
	mem[1215] = 4'b0000;
	mem[1216] = 4'b0000;
	mem[1217] = 4'b0001;
	mem[1218] = 4'b0000;
	mem[1219] = 4'b0000;
	mem[1220] = 4'b0000;
	mem[1221] = 4'b0000;
	mem[1222] = 4'b0000;
	mem[1223] = 4'b1100;
	mem[1224] = 4'b1111;
	mem[1225] = 4'b1111;
	mem[1226] = 4'b1111;
	mem[1227] = 4'b1111;
	mem[1228] = 4'b1111;
	mem[1229] = 4'b1111;
	mem[1230] = 4'b1111;
	mem[1231] = 4'b1111;
	mem[1232] = 4'b1111;
	mem[1233] = 4'b1111;
	mem[1234] = 4'b1111;
	mem[1235] = 4'b1111;
	mem[1236] = 4'b1111;
	mem[1237] = 4'b1111;
	mem[1238] = 4'b1111;
	mem[1239] = 4'b1111;
	mem[1240] = 4'b1111;
	mem[1241] = 4'b1111;
	mem[1242] = 4'b1111;
	mem[1243] = 4'b1111;
	mem[1244] = 4'b1111;
	mem[1245] = 4'b1111;
	mem[1246] = 4'b1111;
	mem[1247] = 4'b1111;
	mem[1248] = 4'b1111;
	mem[1249] = 4'b1111;
	mem[1250] = 4'b1111;
	mem[1251] = 4'b1101;
	mem[1252] = 4'b1110;
	mem[1253] = 4'b1111;
	mem[1254] = 4'b1111;
	mem[1255] = 4'b1101;
	mem[1256] = 4'b1101;
	mem[1257] = 4'b0101;
	mem[1258] = 4'b0000;
	mem[1259] = 4'b0000;
	mem[1260] = 4'b0000;
	mem[1261] = 4'b0000;
	mem[1262] = 4'b0001;
	mem[1263] = 4'b0001;
	mem[1264] = 4'b0000;
	mem[1265] = 4'b0000;
	mem[1266] = 4'b0000;
	mem[1267] = 4'b0000;
	mem[1268] = 4'b0000;
	mem[1269] = 4'b0000;
	mem[1270] = 4'b0000;
	mem[1271] = 4'b0000;
	mem[1272] = 4'b0000;
	mem[1273] = 4'b0000;
	mem[1274] = 4'b0000;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0111;
	mem[1284] = 4'b1100;
	mem[1285] = 4'b1101;
	mem[1286] = 4'b1110;
	mem[1287] = 4'b1110;
	mem[1288] = 4'b1110;
	mem[1289] = 4'b1110;
	mem[1290] = 4'b1110;
	mem[1291] = 4'b1101;
	mem[1292] = 4'b1100;
	mem[1293] = 4'b1100;
	mem[1294] = 4'b1100;
	mem[1295] = 4'b1100;
	mem[1296] = 4'b1100;
	mem[1297] = 4'b1100;
	mem[1298] = 4'b1100;
	mem[1299] = 4'b1100;
	mem[1300] = 4'b1111;
	mem[1301] = 4'b1111;
	mem[1302] = 4'b1111;
	mem[1303] = 4'b1111;
	mem[1304] = 4'b1111;
	mem[1305] = 4'b1111;
	mem[1306] = 4'b1111;
	mem[1307] = 4'b1111;
	mem[1308] = 4'b1111;
	mem[1309] = 4'b1111;
	mem[1310] = 4'b1111;
	mem[1311] = 4'b1111;
	mem[1312] = 4'b1111;
	mem[1313] = 4'b1111;
	mem[1314] = 4'b1111;
	mem[1315] = 4'b1111;
	mem[1316] = 4'b1111;
	mem[1317] = 4'b0100;
	mem[1318] = 4'b0000;
	mem[1319] = 4'b0000;
	mem[1320] = 4'b0000;
	mem[1321] = 4'b0000;
	mem[1322] = 4'b0000;
	mem[1323] = 4'b0000;
	mem[1324] = 4'b0000;
	mem[1325] = 4'b0000;
	mem[1326] = 4'b0000;
	mem[1327] = 4'b0000;
	mem[1328] = 4'b0000;
	mem[1329] = 4'b0000;
	mem[1330] = 4'b0000;
	mem[1331] = 4'b0000;
	mem[1332] = 4'b0000;
	mem[1333] = 4'b0000;
	mem[1334] = 4'b0000;
	mem[1335] = 4'b0000;
	mem[1336] = 4'b0000;
	mem[1337] = 4'b0001;
	mem[1338] = 4'b0001;
	mem[1339] = 4'b0000;
	mem[1340] = 4'b0000;
	mem[1341] = 4'b0000;
	mem[1342] = 4'b0000;
	mem[1343] = 4'b0000;
	mem[1344] = 4'b0000;
	mem[1345] = 4'b0001;
	mem[1346] = 4'b0000;
	mem[1347] = 4'b0000;
	mem[1348] = 4'b0000;
	mem[1349] = 4'b0000;
	mem[1350] = 4'b0000;
	mem[1351] = 4'b1100;
	mem[1352] = 4'b1111;
	mem[1353] = 4'b1111;
	mem[1354] = 4'b1111;
	mem[1355] = 4'b1111;
	mem[1356] = 4'b1111;
	mem[1357] = 4'b1111;
	mem[1358] = 4'b1111;
	mem[1359] = 4'b1111;
	mem[1360] = 4'b1111;
	mem[1361] = 4'b1111;
	mem[1362] = 4'b1111;
	mem[1363] = 4'b1111;
	mem[1364] = 4'b1111;
	mem[1365] = 4'b1111;
	mem[1366] = 4'b1111;
	mem[1367] = 4'b1111;
	mem[1368] = 4'b1111;
	mem[1369] = 4'b1111;
	mem[1370] = 4'b1111;
	mem[1371] = 4'b1111;
	mem[1372] = 4'b1111;
	mem[1373] = 4'b1111;
	mem[1374] = 4'b1111;
	mem[1375] = 4'b1111;
	mem[1376] = 4'b1111;
	mem[1377] = 4'b1111;
	mem[1378] = 4'b1110;
	mem[1379] = 4'b1101;
	mem[1380] = 4'b1111;
	mem[1381] = 4'b1111;
	mem[1382] = 4'b1110;
	mem[1383] = 4'b1110;
	mem[1384] = 4'b1110;
	mem[1385] = 4'b0101;
	mem[1386] = 4'b0000;
	mem[1387] = 4'b0000;
	mem[1388] = 4'b0000;
	mem[1389] = 4'b0000;
	mem[1390] = 4'b0000;
	mem[1391] = 4'b0000;
	mem[1392] = 4'b0000;
	mem[1393] = 4'b0000;
	mem[1394] = 4'b0000;
	mem[1395] = 4'b0000;
	mem[1396] = 4'b0000;
	mem[1397] = 4'b0000;
	mem[1398] = 4'b0000;
	mem[1399] = 4'b0000;
	mem[1400] = 4'b0000;
	mem[1401] = 4'b0000;
	mem[1402] = 4'b0000;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0111;
	mem[1412] = 4'b1100;
	mem[1413] = 4'b1101;
	mem[1414] = 4'b1110;
	mem[1415] = 4'b1110;
	mem[1416] = 4'b1110;
	mem[1417] = 4'b1101;
	mem[1418] = 4'b1100;
	mem[1419] = 4'b1100;
	mem[1420] = 4'b1100;
	mem[1421] = 4'b1100;
	mem[1422] = 4'b1100;
	mem[1423] = 4'b1100;
	mem[1424] = 4'b1100;
	mem[1425] = 4'b1100;
	mem[1426] = 4'b1100;
	mem[1427] = 4'b1100;
	mem[1428] = 4'b1111;
	mem[1429] = 4'b1111;
	mem[1430] = 4'b1111;
	mem[1431] = 4'b1111;
	mem[1432] = 4'b1111;
	mem[1433] = 4'b1111;
	mem[1434] = 4'b1111;
	mem[1435] = 4'b1111;
	mem[1436] = 4'b1111;
	mem[1437] = 4'b1111;
	mem[1438] = 4'b1111;
	mem[1439] = 4'b1111;
	mem[1440] = 4'b1111;
	mem[1441] = 4'b1111;
	mem[1442] = 4'b1111;
	mem[1443] = 4'b1111;
	mem[1444] = 4'b1111;
	mem[1445] = 4'b0100;
	mem[1446] = 4'b0000;
	mem[1447] = 4'b0000;
	mem[1448] = 4'b0000;
	mem[1449] = 4'b0000;
	mem[1450] = 4'b0000;
	mem[1451] = 4'b0000;
	mem[1452] = 4'b0000;
	mem[1453] = 4'b0000;
	mem[1454] = 4'b0000;
	mem[1455] = 4'b0000;
	mem[1456] = 4'b0000;
	mem[1457] = 4'b0000;
	mem[1458] = 4'b0000;
	mem[1459] = 4'b0000;
	mem[1460] = 4'b0000;
	mem[1461] = 4'b0000;
	mem[1462] = 4'b0000;
	mem[1463] = 4'b0001;
	mem[1464] = 4'b0001;
	mem[1465] = 4'b0000;
	mem[1466] = 4'b0000;
	mem[1467] = 4'b0000;
	mem[1468] = 4'b0000;
	mem[1469] = 4'b0000;
	mem[1470] = 4'b0000;
	mem[1471] = 4'b0000;
	mem[1472] = 4'b0001;
	mem[1473] = 4'b0001;
	mem[1474] = 4'b0000;
	mem[1475] = 4'b0000;
	mem[1476] = 4'b0000;
	mem[1477] = 4'b0000;
	mem[1478] = 4'b0000;
	mem[1479] = 4'b1100;
	mem[1480] = 4'b1111;
	mem[1481] = 4'b1111;
	mem[1482] = 4'b1111;
	mem[1483] = 4'b1111;
	mem[1484] = 4'b1111;
	mem[1485] = 4'b1111;
	mem[1486] = 4'b1111;
	mem[1487] = 4'b1111;
	mem[1488] = 4'b1111;
	mem[1489] = 4'b1111;
	mem[1490] = 4'b1111;
	mem[1491] = 4'b1111;
	mem[1492] = 4'b1111;
	mem[1493] = 4'b1111;
	mem[1494] = 4'b1111;
	mem[1495] = 4'b1111;
	mem[1496] = 4'b1111;
	mem[1497] = 4'b1111;
	mem[1498] = 4'b1111;
	mem[1499] = 4'b1111;
	mem[1500] = 4'b1111;
	mem[1501] = 4'b1111;
	mem[1502] = 4'b1111;
	mem[1503] = 4'b1111;
	mem[1504] = 4'b1111;
	mem[1505] = 4'b1111;
	mem[1506] = 4'b1111;
	mem[1507] = 4'b1110;
	mem[1508] = 4'b1111;
	mem[1509] = 4'b1111;
	mem[1510] = 4'b1101;
	mem[1511] = 4'b1111;
	mem[1512] = 4'b1111;
	mem[1513] = 4'b0101;
	mem[1514] = 4'b0000;
	mem[1515] = 4'b0000;
	mem[1516] = 4'b0001;
	mem[1517] = 4'b0000;
	mem[1518] = 4'b0000;
	mem[1519] = 4'b0000;
	mem[1520] = 4'b0000;
	mem[1521] = 4'b0000;
	mem[1522] = 4'b0000;
	mem[1523] = 4'b0000;
	mem[1524] = 4'b0000;
	mem[1525] = 4'b0000;
	mem[1526] = 4'b0000;
	mem[1527] = 4'b0000;
	mem[1528] = 4'b0000;
	mem[1529] = 4'b0000;
	mem[1530] = 4'b0000;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0001;
	mem[1540] = 4'b0001;
	mem[1541] = 4'b0101;
	mem[1542] = 4'b1000;
	mem[1543] = 4'b1000;
	mem[1544] = 4'b0101;
	mem[1545] = 4'b0001;
	mem[1546] = 4'b0001;
	mem[1547] = 4'b0001;
	mem[1548] = 4'b0001;
	mem[1549] = 4'b0001;
	mem[1550] = 4'b0001;
	mem[1551] = 4'b0001;
	mem[1552] = 4'b0001;
	mem[1553] = 4'b0001;
	mem[1554] = 4'b0001;
	mem[1555] = 4'b0001;
	mem[1556] = 4'b0001;
	mem[1557] = 4'b0010;
	mem[1558] = 4'b0010;
	mem[1559] = 4'b0010;
	mem[1560] = 4'b0010;
	mem[1561] = 4'b0010;
	mem[1562] = 4'b0010;
	mem[1563] = 4'b0010;
	mem[1564] = 4'b0010;
	mem[1565] = 4'b0010;
	mem[1566] = 4'b0010;
	mem[1567] = 4'b0010;
	mem[1568] = 4'b0010;
	mem[1569] = 4'b0010;
	mem[1570] = 4'b0010;
	mem[1571] = 4'b0010;
	mem[1572] = 4'b0010;
	mem[1573] = 4'b1011;
	mem[1574] = 4'b1101;
	mem[1575] = 4'b1101;
	mem[1576] = 4'b1101;
	mem[1577] = 4'b1101;
	mem[1578] = 4'b1101;
	mem[1579] = 4'b1100;
	mem[1580] = 4'b1100;
	mem[1581] = 4'b1100;
	mem[1582] = 4'b1100;
	mem[1583] = 4'b1101;
	mem[1584] = 4'b1101;
	mem[1585] = 4'b1101;
	mem[1586] = 4'b1101;
	mem[1587] = 4'b1110;
	mem[1588] = 4'b1101;
	mem[1589] = 4'b1101;
	mem[1590] = 4'b0110;
	mem[1591] = 4'b0000;
	mem[1592] = 4'b0000;
	mem[1593] = 4'b0000;
	mem[1594] = 4'b0000;
	mem[1595] = 4'b0000;
	mem[1596] = 4'b0000;
	mem[1597] = 4'b0000;
	mem[1598] = 4'b0000;
	mem[1599] = 4'b0000;
	mem[1600] = 4'b0001;
	mem[1601] = 4'b0000;
	mem[1602] = 4'b0000;
	mem[1603] = 4'b0000;
	mem[1604] = 4'b0000;
	mem[1605] = 4'b0000;
	mem[1606] = 4'b0000;
	mem[1607] = 4'b0001;
	mem[1608] = 4'b0010;
	mem[1609] = 4'b0010;
	mem[1610] = 4'b0010;
	mem[1611] = 4'b0010;
	mem[1612] = 4'b0010;
	mem[1613] = 4'b0010;
	mem[1614] = 4'b0010;
	mem[1615] = 4'b0010;
	mem[1616] = 4'b0010;
	mem[1617] = 4'b0010;
	mem[1618] = 4'b0010;
	mem[1619] = 4'b0010;
	mem[1620] = 4'b0010;
	mem[1621] = 4'b0010;
	mem[1622] = 4'b0010;
	mem[1623] = 4'b0010;
	mem[1624] = 4'b0010;
	mem[1625] = 4'b0010;
	mem[1626] = 4'b0010;
	mem[1627] = 4'b0010;
	mem[1628] = 4'b0010;
	mem[1629] = 4'b0010;
	mem[1630] = 4'b0010;
	mem[1631] = 4'b0010;
	mem[1632] = 4'b0010;
	mem[1633] = 4'b0010;
	mem[1634] = 4'b0010;
	mem[1635] = 4'b0011;
	mem[1636] = 4'b0010;
	mem[1637] = 4'b0010;
	mem[1638] = 4'b0010;
	mem[1639] = 4'b0011;
	mem[1640] = 4'b0010;
	mem[1641] = 4'b0111;
	mem[1642] = 4'b1010;
	mem[1643] = 4'b1010;
	mem[1644] = 4'b1011;
	mem[1645] = 4'b1011;
	mem[1646] = 4'b1011;
	mem[1647] = 4'b1011;
	mem[1648] = 4'b1011;
	mem[1649] = 4'b1011;
	mem[1650] = 4'b1011;
	mem[1651] = 4'b1011;
	mem[1652] = 4'b1011;
	mem[1653] = 4'b1011;
	mem[1654] = 4'b1011;
	mem[1655] = 4'b1011;
	mem[1656] = 4'b1011;
	mem[1657] = 4'b1010;
	mem[1658] = 4'b0010;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0000;
	mem[1668] = 4'b0000;
	mem[1669] = 4'b0100;
	mem[1670] = 4'b0111;
	mem[1671] = 4'b0011;
	mem[1672] = 4'b0000;
	mem[1673] = 4'b0000;
	mem[1674] = 4'b0000;
	mem[1675] = 4'b0000;
	mem[1676] = 4'b0000;
	mem[1677] = 4'b0000;
	mem[1678] = 4'b0000;
	mem[1679] = 4'b0000;
	mem[1680] = 4'b0000;
	mem[1681] = 4'b0000;
	mem[1682] = 4'b0000;
	mem[1683] = 4'b0000;
	mem[1684] = 4'b0000;
	mem[1685] = 4'b0000;
	mem[1686] = 4'b0000;
	mem[1687] = 4'b0000;
	mem[1688] = 4'b0000;
	mem[1689] = 4'b0000;
	mem[1690] = 4'b0000;
	mem[1691] = 4'b0000;
	mem[1692] = 4'b0000;
	mem[1693] = 4'b0000;
	mem[1694] = 4'b0000;
	mem[1695] = 4'b0000;
	mem[1696] = 4'b0000;
	mem[1697] = 4'b0000;
	mem[1698] = 4'b0000;
	mem[1699] = 4'b0000;
	mem[1700] = 4'b0000;
	mem[1701] = 4'b1100;
	mem[1702] = 4'b1111;
	mem[1703] = 4'b1111;
	mem[1704] = 4'b1111;
	mem[1705] = 4'b1110;
	mem[1706] = 4'b1101;
	mem[1707] = 4'b1101;
	mem[1708] = 4'b1101;
	mem[1709] = 4'b1101;
	mem[1710] = 4'b1101;
	mem[1711] = 4'b1101;
	mem[1712] = 4'b1111;
	mem[1713] = 4'b1111;
	mem[1714] = 4'b1111;
	mem[1715] = 4'b1111;
	mem[1716] = 4'b1111;
	mem[1717] = 4'b1111;
	mem[1718] = 4'b0110;
	mem[1719] = 4'b0000;
	mem[1720] = 4'b0000;
	mem[1721] = 4'b0000;
	mem[1722] = 4'b0000;
	mem[1723] = 4'b0000;
	mem[1724] = 4'b0000;
	mem[1725] = 4'b0000;
	mem[1726] = 4'b0000;
	mem[1727] = 4'b0001;
	mem[1728] = 4'b0001;
	mem[1729] = 4'b0000;
	mem[1730] = 4'b0000;
	mem[1731] = 4'b0000;
	mem[1732] = 4'b0000;
	mem[1733] = 4'b0000;
	mem[1734] = 4'b0000;
	mem[1735] = 4'b0000;
	mem[1736] = 4'b0000;
	mem[1737] = 4'b0000;
	mem[1738] = 4'b0000;
	mem[1739] = 4'b0000;
	mem[1740] = 4'b0000;
	mem[1741] = 4'b0000;
	mem[1742] = 4'b0000;
	mem[1743] = 4'b0000;
	mem[1744] = 4'b0000;
	mem[1745] = 4'b0000;
	mem[1746] = 4'b0000;
	mem[1747] = 4'b0000;
	mem[1748] = 4'b0000;
	mem[1749] = 4'b0000;
	mem[1750] = 4'b0000;
	mem[1751] = 4'b0000;
	mem[1752] = 4'b0000;
	mem[1753] = 4'b0000;
	mem[1754] = 4'b0000;
	mem[1755] = 4'b0000;
	mem[1756] = 4'b0000;
	mem[1757] = 4'b0000;
	mem[1758] = 4'b0000;
	mem[1759] = 4'b0000;
	mem[1760] = 4'b0000;
	mem[1761] = 4'b0000;
	mem[1762] = 4'b0000;
	mem[1763] = 4'b0000;
	mem[1764] = 4'b0000;
	mem[1765] = 4'b0000;
	mem[1766] = 4'b0000;
	mem[1767] = 4'b0000;
	mem[1768] = 4'b0000;
	mem[1769] = 4'b0111;
	mem[1770] = 4'b1100;
	mem[1771] = 4'b1100;
	mem[1772] = 4'b1100;
	mem[1773] = 4'b1100;
	mem[1774] = 4'b1100;
	mem[1775] = 4'b1100;
	mem[1776] = 4'b1100;
	mem[1777] = 4'b1100;
	mem[1778] = 4'b1100;
	mem[1779] = 4'b1100;
	mem[1780] = 4'b1100;
	mem[1781] = 4'b1100;
	mem[1782] = 4'b1100;
	mem[1783] = 4'b1100;
	mem[1784] = 4'b1100;
	mem[1785] = 4'b1100;
	mem[1786] = 4'b0010;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0000;
	mem[1796] = 4'b0000;
	mem[1797] = 4'b0100;
	mem[1798] = 4'b0011;
	mem[1799] = 4'b0000;
	mem[1800] = 4'b0000;
	mem[1801] = 4'b0000;
	mem[1802] = 4'b0000;
	mem[1803] = 4'b0000;
	mem[1804] = 4'b0000;
	mem[1805] = 4'b0000;
	mem[1806] = 4'b0000;
	mem[1807] = 4'b0000;
	mem[1808] = 4'b0000;
	mem[1809] = 4'b0000;
	mem[1810] = 4'b0000;
	mem[1811] = 4'b0000;
	mem[1812] = 4'b0000;
	mem[1813] = 4'b0000;
	mem[1814] = 4'b0000;
	mem[1815] = 4'b0000;
	mem[1816] = 4'b0000;
	mem[1817] = 4'b0000;
	mem[1818] = 4'b0000;
	mem[1819] = 4'b0000;
	mem[1820] = 4'b0000;
	mem[1821] = 4'b0000;
	mem[1822] = 4'b0000;
	mem[1823] = 4'b0000;
	mem[1824] = 4'b0000;
	mem[1825] = 4'b0000;
	mem[1826] = 4'b0000;
	mem[1827] = 4'b0000;
	mem[1828] = 4'b0000;
	mem[1829] = 4'b1100;
	mem[1830] = 4'b1111;
	mem[1831] = 4'b1111;
	mem[1832] = 4'b1110;
	mem[1833] = 4'b1101;
	mem[1834] = 4'b1101;
	mem[1835] = 4'b1101;
	mem[1836] = 4'b1101;
	mem[1837] = 4'b1101;
	mem[1838] = 4'b1101;
	mem[1839] = 4'b1101;
	mem[1840] = 4'b1101;
	mem[1841] = 4'b1111;
	mem[1842] = 4'b1111;
	mem[1843] = 4'b1111;
	mem[1844] = 4'b1111;
	mem[1845] = 4'b1111;
	mem[1846] = 4'b0110;
	mem[1847] = 4'b0000;
	mem[1848] = 4'b0000;
	mem[1849] = 4'b0000;
	mem[1850] = 4'b0000;
	mem[1851] = 4'b0000;
	mem[1852] = 4'b0000;
	mem[1853] = 4'b0000;
	mem[1854] = 4'b0001;
	mem[1855] = 4'b0001;
	mem[1856] = 4'b0000;
	mem[1857] = 4'b0000;
	mem[1858] = 4'b0000;
	mem[1859] = 4'b0000;
	mem[1860] = 4'b0000;
	mem[1861] = 4'b0000;
	mem[1862] = 4'b0000;
	mem[1863] = 4'b0000;
	mem[1864] = 4'b0000;
	mem[1865] = 4'b0000;
	mem[1866] = 4'b0000;
	mem[1867] = 4'b0000;
	mem[1868] = 4'b0000;
	mem[1869] = 4'b0000;
	mem[1870] = 4'b0000;
	mem[1871] = 4'b0000;
	mem[1872] = 4'b0000;
	mem[1873] = 4'b0000;
	mem[1874] = 4'b0000;
	mem[1875] = 4'b0000;
	mem[1876] = 4'b0000;
	mem[1877] = 4'b0000;
	mem[1878] = 4'b0000;
	mem[1879] = 4'b0000;
	mem[1880] = 4'b0000;
	mem[1881] = 4'b0000;
	mem[1882] = 4'b0000;
	mem[1883] = 4'b0000;
	mem[1884] = 4'b0000;
	mem[1885] = 4'b0000;
	mem[1886] = 4'b0000;
	mem[1887] = 4'b0000;
	mem[1888] = 4'b0000;
	mem[1889] = 4'b0000;
	mem[1890] = 4'b0000;
	mem[1891] = 4'b0000;
	mem[1892] = 4'b0000;
	mem[1893] = 4'b0000;
	mem[1894] = 4'b0000;
	mem[1895] = 4'b0000;
	mem[1896] = 4'b0000;
	mem[1897] = 4'b0111;
	mem[1898] = 4'b1101;
	mem[1899] = 4'b1100;
	mem[1900] = 4'b1100;
	mem[1901] = 4'b1100;
	mem[1902] = 4'b1100;
	mem[1903] = 4'b1100;
	mem[1904] = 4'b1100;
	mem[1905] = 4'b1100;
	mem[1906] = 4'b1100;
	mem[1907] = 4'b1100;
	mem[1908] = 4'b1100;
	mem[1909] = 4'b1100;
	mem[1910] = 4'b1100;
	mem[1911] = 4'b1100;
	mem[1912] = 4'b1100;
	mem[1913] = 4'b1100;
	mem[1914] = 4'b0010;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0000;
	mem[1924] = 4'b0000;
	mem[1925] = 4'b0000;
	mem[1926] = 4'b0000;
	mem[1927] = 4'b0000;
	mem[1928] = 4'b0000;
	mem[1929] = 4'b0000;
	mem[1930] = 4'b0000;
	mem[1931] = 4'b0000;
	mem[1932] = 4'b0000;
	mem[1933] = 4'b0000;
	mem[1934] = 4'b0000;
	mem[1935] = 4'b0000;
	mem[1936] = 4'b0000;
	mem[1937] = 4'b0000;
	mem[1938] = 4'b0000;
	mem[1939] = 4'b0000;
	mem[1940] = 4'b0000;
	mem[1941] = 4'b0000;
	mem[1942] = 4'b0000;
	mem[1943] = 4'b0000;
	mem[1944] = 4'b0000;
	mem[1945] = 4'b0000;
	mem[1946] = 4'b0000;
	mem[1947] = 4'b0000;
	mem[1948] = 4'b0000;
	mem[1949] = 4'b0000;
	mem[1950] = 4'b0000;
	mem[1951] = 4'b0000;
	mem[1952] = 4'b0000;
	mem[1953] = 4'b0000;
	mem[1954] = 4'b0000;
	mem[1955] = 4'b0000;
	mem[1956] = 4'b0000;
	mem[1957] = 4'b1100;
	mem[1958] = 4'b1111;
	mem[1959] = 4'b1111;
	mem[1960] = 4'b1101;
	mem[1961] = 4'b1101;
	mem[1962] = 4'b1101;
	mem[1963] = 4'b1101;
	mem[1964] = 4'b1101;
	mem[1965] = 4'b1101;
	mem[1966] = 4'b1101;
	mem[1967] = 4'b1101;
	mem[1968] = 4'b1101;
	mem[1969] = 4'b1101;
	mem[1970] = 4'b1111;
	mem[1971] = 4'b1111;
	mem[1972] = 4'b1111;
	mem[1973] = 4'b1111;
	mem[1974] = 4'b0101;
	mem[1975] = 4'b0000;
	mem[1976] = 4'b0000;
	mem[1977] = 4'b0000;
	mem[1978] = 4'b0000;
	mem[1979] = 4'b0000;
	mem[1980] = 4'b0000;
	mem[1981] = 4'b0001;
	mem[1982] = 4'b0001;
	mem[1983] = 4'b0000;
	mem[1984] = 4'b0000;
	mem[1985] = 4'b0000;
	mem[1986] = 4'b0000;
	mem[1987] = 4'b0000;
	mem[1988] = 4'b0000;
	mem[1989] = 4'b0000;
	mem[1990] = 4'b0000;
	mem[1991] = 4'b0000;
	mem[1992] = 4'b0000;
	mem[1993] = 4'b0000;
	mem[1994] = 4'b0000;
	mem[1995] = 4'b0000;
	mem[1996] = 4'b0000;
	mem[1997] = 4'b0000;
	mem[1998] = 4'b0000;
	mem[1999] = 4'b0000;
	mem[2000] = 4'b0000;
	mem[2001] = 4'b0000;
	mem[2002] = 4'b0000;
	mem[2003] = 4'b0000;
	mem[2004] = 4'b0000;
	mem[2005] = 4'b0000;
	mem[2006] = 4'b0000;
	mem[2007] = 4'b0000;
	mem[2008] = 4'b0000;
	mem[2009] = 4'b0000;
	mem[2010] = 4'b0000;
	mem[2011] = 4'b0000;
	mem[2012] = 4'b0000;
	mem[2013] = 4'b0000;
	mem[2014] = 4'b0000;
	mem[2015] = 4'b0000;
	mem[2016] = 4'b0000;
	mem[2017] = 4'b0000;
	mem[2018] = 4'b0000;
	mem[2019] = 4'b0000;
	mem[2020] = 4'b0000;
	mem[2021] = 4'b0000;
	mem[2022] = 4'b0000;
	mem[2023] = 4'b0000;
	mem[2024] = 4'b0001;
	mem[2025] = 4'b1000;
	mem[2026] = 4'b1100;
	mem[2027] = 4'b1100;
	mem[2028] = 4'b1100;
	mem[2029] = 4'b1100;
	mem[2030] = 4'b1100;
	mem[2031] = 4'b1100;
	mem[2032] = 4'b1100;
	mem[2033] = 4'b1100;
	mem[2034] = 4'b1100;
	mem[2035] = 4'b1100;
	mem[2036] = 4'b1100;
	mem[2037] = 4'b1100;
	mem[2038] = 4'b1100;
	mem[2039] = 4'b1100;
	mem[2040] = 4'b1100;
	mem[2041] = 4'b1100;
	mem[2042] = 4'b0010;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0000;
	mem[2052] = 4'b0000;
	mem[2053] = 4'b0000;
	mem[2054] = 4'b0000;
	mem[2055] = 4'b0000;
	mem[2056] = 4'b0000;
	mem[2057] = 4'b0000;
	mem[2058] = 4'b0000;
	mem[2059] = 4'b0000;
	mem[2060] = 4'b0000;
	mem[2061] = 4'b0000;
	mem[2062] = 4'b0000;
	mem[2063] = 4'b0000;
	mem[2064] = 4'b0000;
	mem[2065] = 4'b0000;
	mem[2066] = 4'b0000;
	mem[2067] = 4'b0000;
	mem[2068] = 4'b0000;
	mem[2069] = 4'b0000;
	mem[2070] = 4'b0000;
	mem[2071] = 4'b0000;
	mem[2072] = 4'b0000;
	mem[2073] = 4'b0000;
	mem[2074] = 4'b0000;
	mem[2075] = 4'b0000;
	mem[2076] = 4'b0000;
	mem[2077] = 4'b0000;
	mem[2078] = 4'b0000;
	mem[2079] = 4'b0000;
	mem[2080] = 4'b0000;
	mem[2081] = 4'b0000;
	mem[2082] = 4'b0000;
	mem[2083] = 4'b0000;
	mem[2084] = 4'b0000;
	mem[2085] = 4'b1100;
	mem[2086] = 4'b1111;
	mem[2087] = 4'b1111;
	mem[2088] = 4'b1101;
	mem[2089] = 4'b1101;
	mem[2090] = 4'b1110;
	mem[2091] = 4'b1111;
	mem[2092] = 4'b1111;
	mem[2093] = 4'b1111;
	mem[2094] = 4'b1101;
	mem[2095] = 4'b1101;
	mem[2096] = 4'b1101;
	mem[2097] = 4'b1101;
	mem[2098] = 4'b1101;
	mem[2099] = 4'b1111;
	mem[2100] = 4'b1111;
	mem[2101] = 4'b1111;
	mem[2102] = 4'b0110;
	mem[2103] = 4'b0001;
	mem[2104] = 4'b0001;
	mem[2105] = 4'b0000;
	mem[2106] = 4'b0001;
	mem[2107] = 4'b0001;
	mem[2108] = 4'b0001;
	mem[2109] = 4'b0000;
	mem[2110] = 4'b0000;
	mem[2111] = 4'b0000;
	mem[2112] = 4'b0000;
	mem[2113] = 4'b0000;
	mem[2114] = 4'b0000;
	mem[2115] = 4'b0000;
	mem[2116] = 4'b0000;
	mem[2117] = 4'b0000;
	mem[2118] = 4'b0000;
	mem[2119] = 4'b0000;
	mem[2120] = 4'b0000;
	mem[2121] = 4'b0000;
	mem[2122] = 4'b0000;
	mem[2123] = 4'b0000;
	mem[2124] = 4'b0000;
	mem[2125] = 4'b0000;
	mem[2126] = 4'b0000;
	mem[2127] = 4'b0000;
	mem[2128] = 4'b0000;
	mem[2129] = 4'b0000;
	mem[2130] = 4'b0000;
	mem[2131] = 4'b0000;
	mem[2132] = 4'b0000;
	mem[2133] = 4'b0000;
	mem[2134] = 4'b0000;
	mem[2135] = 4'b0000;
	mem[2136] = 4'b0000;
	mem[2137] = 4'b0000;
	mem[2138] = 4'b0000;
	mem[2139] = 4'b0000;
	mem[2140] = 4'b0000;
	mem[2141] = 4'b0000;
	mem[2142] = 4'b0000;
	mem[2143] = 4'b0000;
	mem[2144] = 4'b0000;
	mem[2145] = 4'b0000;
	mem[2146] = 4'b0000;
	mem[2147] = 4'b0000;
	mem[2148] = 4'b0000;
	mem[2149] = 4'b0000;
	mem[2150] = 4'b0000;
	mem[2151] = 4'b0001;
	mem[2152] = 4'b0001;
	mem[2153] = 4'b1000;
	mem[2154] = 4'b1100;
	mem[2155] = 4'b1100;
	mem[2156] = 4'b1100;
	mem[2157] = 4'b1100;
	mem[2158] = 4'b1100;
	mem[2159] = 4'b1100;
	mem[2160] = 4'b1100;
	mem[2161] = 4'b1100;
	mem[2162] = 4'b1100;
	mem[2163] = 4'b1100;
	mem[2164] = 4'b1100;
	mem[2165] = 4'b1100;
	mem[2166] = 4'b1100;
	mem[2167] = 4'b1100;
	mem[2168] = 4'b1100;
	mem[2169] = 4'b1100;
	mem[2170] = 4'b0010;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0000;
	mem[2180] = 4'b0000;
	mem[2181] = 4'b0000;
	mem[2182] = 4'b0000;
	mem[2183] = 4'b0000;
	mem[2184] = 4'b0000;
	mem[2185] = 4'b0000;
	mem[2186] = 4'b0000;
	mem[2187] = 4'b0000;
	mem[2188] = 4'b0000;
	mem[2189] = 4'b0000;
	mem[2190] = 4'b0000;
	mem[2191] = 4'b0000;
	mem[2192] = 4'b0000;
	mem[2193] = 4'b0000;
	mem[2194] = 4'b0000;
	mem[2195] = 4'b0000;
	mem[2196] = 4'b0000;
	mem[2197] = 4'b0000;
	mem[2198] = 4'b0000;
	mem[2199] = 4'b0000;
	mem[2200] = 4'b0000;
	mem[2201] = 4'b0000;
	mem[2202] = 4'b0000;
	mem[2203] = 4'b0000;
	mem[2204] = 4'b0000;
	mem[2205] = 4'b0000;
	mem[2206] = 4'b0000;
	mem[2207] = 4'b0000;
	mem[2208] = 4'b0000;
	mem[2209] = 4'b0000;
	mem[2210] = 4'b0000;
	mem[2211] = 4'b0000;
	mem[2212] = 4'b0000;
	mem[2213] = 4'b1011;
	mem[2214] = 4'b1111;
	mem[2215] = 4'b1111;
	mem[2216] = 4'b1101;
	mem[2217] = 4'b1110;
	mem[2218] = 4'b1111;
	mem[2219] = 4'b1111;
	mem[2220] = 4'b1111;
	mem[2221] = 4'b1111;
	mem[2222] = 4'b1111;
	mem[2223] = 4'b1101;
	mem[2224] = 4'b1101;
	mem[2225] = 4'b1101;
	mem[2226] = 4'b1101;
	mem[2227] = 4'b1101;
	mem[2228] = 4'b1111;
	mem[2229] = 4'b1111;
	mem[2230] = 4'b0110;
	mem[2231] = 4'b0000;
	mem[2232] = 4'b0000;
	mem[2233] = 4'b0000;
	mem[2234] = 4'b0000;
	mem[2235] = 4'b0000;
	mem[2236] = 4'b0000;
	mem[2237] = 4'b0000;
	mem[2238] = 4'b0000;
	mem[2239] = 4'b0000;
	mem[2240] = 4'b0000;
	mem[2241] = 4'b0000;
	mem[2242] = 4'b0000;
	mem[2243] = 4'b0000;
	mem[2244] = 4'b0000;
	mem[2245] = 4'b0000;
	mem[2246] = 4'b0000;
	mem[2247] = 4'b0000;
	mem[2248] = 4'b0000;
	mem[2249] = 4'b0000;
	mem[2250] = 4'b0000;
	mem[2251] = 4'b0000;
	mem[2252] = 4'b0000;
	mem[2253] = 4'b0000;
	mem[2254] = 4'b0000;
	mem[2255] = 4'b0000;
	mem[2256] = 4'b0000;
	mem[2257] = 4'b0000;
	mem[2258] = 4'b0000;
	mem[2259] = 4'b0000;
	mem[2260] = 4'b0000;
	mem[2261] = 4'b0000;
	mem[2262] = 4'b0000;
	mem[2263] = 4'b0000;
	mem[2264] = 4'b0000;
	mem[2265] = 4'b0000;
	mem[2266] = 4'b0000;
	mem[2267] = 4'b0000;
	mem[2268] = 4'b0000;
	mem[2269] = 4'b0000;
	mem[2270] = 4'b0000;
	mem[2271] = 4'b0000;
	mem[2272] = 4'b0000;
	mem[2273] = 4'b0000;
	mem[2274] = 4'b0000;
	mem[2275] = 4'b0000;
	mem[2276] = 4'b0000;
	mem[2277] = 4'b0000;
	mem[2278] = 4'b0000;
	mem[2279] = 4'b0000;
	mem[2280] = 4'b0000;
	mem[2281] = 4'b1000;
	mem[2282] = 4'b1100;
	mem[2283] = 4'b1100;
	mem[2284] = 4'b1100;
	mem[2285] = 4'b1100;
	mem[2286] = 4'b1100;
	mem[2287] = 4'b1100;
	mem[2288] = 4'b1100;
	mem[2289] = 4'b1100;
	mem[2290] = 4'b1100;
	mem[2291] = 4'b1100;
	mem[2292] = 4'b1100;
	mem[2293] = 4'b1100;
	mem[2294] = 4'b1100;
	mem[2295] = 4'b1100;
	mem[2296] = 4'b1100;
	mem[2297] = 4'b1100;
	mem[2298] = 4'b0010;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0000;
	mem[2308] = 4'b0000;
	mem[2309] = 4'b0000;
	mem[2310] = 4'b0000;
	mem[2311] = 4'b0000;
	mem[2312] = 4'b0000;
	mem[2313] = 4'b0000;
	mem[2314] = 4'b0000;
	mem[2315] = 4'b0000;
	mem[2316] = 4'b0000;
	mem[2317] = 4'b0000;
	mem[2318] = 4'b0000;
	mem[2319] = 4'b0000;
	mem[2320] = 4'b0000;
	mem[2321] = 4'b0000;
	mem[2322] = 4'b0000;
	mem[2323] = 4'b0000;
	mem[2324] = 4'b0000;
	mem[2325] = 4'b0000;
	mem[2326] = 4'b0000;
	mem[2327] = 4'b0000;
	mem[2328] = 4'b0000;
	mem[2329] = 4'b0000;
	mem[2330] = 4'b0000;
	mem[2331] = 4'b0000;
	mem[2332] = 4'b0000;
	mem[2333] = 4'b0000;
	mem[2334] = 4'b0000;
	mem[2335] = 4'b0000;
	mem[2336] = 4'b0000;
	mem[2337] = 4'b0000;
	mem[2338] = 4'b0000;
	mem[2339] = 4'b0000;
	mem[2340] = 4'b0000;
	mem[2341] = 4'b1010;
	mem[2342] = 4'b1110;
	mem[2343] = 4'b1110;
	mem[2344] = 4'b1101;
	mem[2345] = 4'b1111;
	mem[2346] = 4'b1111;
	mem[2347] = 4'b1111;
	mem[2348] = 4'b1111;
	mem[2349] = 4'b1111;
	mem[2350] = 4'b1111;
	mem[2351] = 4'b1111;
	mem[2352] = 4'b1101;
	mem[2353] = 4'b1101;
	mem[2354] = 4'b1101;
	mem[2355] = 4'b1101;
	mem[2356] = 4'b1101;
	mem[2357] = 4'b1111;
	mem[2358] = 4'b0110;
	mem[2359] = 4'b0000;
	mem[2360] = 4'b0000;
	mem[2361] = 4'b0000;
	mem[2362] = 4'b0000;
	mem[2363] = 4'b0000;
	mem[2364] = 4'b0000;
	mem[2365] = 4'b0000;
	mem[2366] = 4'b0000;
	mem[2367] = 4'b0000;
	mem[2368] = 4'b0000;
	mem[2369] = 4'b0000;
	mem[2370] = 4'b0000;
	mem[2371] = 4'b0000;
	mem[2372] = 4'b0000;
	mem[2373] = 4'b0000;
	mem[2374] = 4'b0000;
	mem[2375] = 4'b0000;
	mem[2376] = 4'b0000;
	mem[2377] = 4'b0000;
	mem[2378] = 4'b0000;
	mem[2379] = 4'b0000;
	mem[2380] = 4'b0000;
	mem[2381] = 4'b0000;
	mem[2382] = 4'b0000;
	mem[2383] = 4'b0000;
	mem[2384] = 4'b0000;
	mem[2385] = 4'b0000;
	mem[2386] = 4'b0000;
	mem[2387] = 4'b0000;
	mem[2388] = 4'b0000;
	mem[2389] = 4'b0000;
	mem[2390] = 4'b0000;
	mem[2391] = 4'b0000;
	mem[2392] = 4'b0000;
	mem[2393] = 4'b0000;
	mem[2394] = 4'b0000;
	mem[2395] = 4'b0000;
	mem[2396] = 4'b0000;
	mem[2397] = 4'b0000;
	mem[2398] = 4'b0000;
	mem[2399] = 4'b0000;
	mem[2400] = 4'b0000;
	mem[2401] = 4'b0000;
	mem[2402] = 4'b0000;
	mem[2403] = 4'b0000;
	mem[2404] = 4'b0000;
	mem[2405] = 4'b0001;
	mem[2406] = 4'b0001;
	mem[2407] = 4'b0000;
	mem[2408] = 4'b0000;
	mem[2409] = 4'b1000;
	mem[2410] = 4'b1100;
	mem[2411] = 4'b1100;
	mem[2412] = 4'b1100;
	mem[2413] = 4'b1100;
	mem[2414] = 4'b1100;
	mem[2415] = 4'b1100;
	mem[2416] = 4'b1100;
	mem[2417] = 4'b1100;
	mem[2418] = 4'b1100;
	mem[2419] = 4'b1100;
	mem[2420] = 4'b1100;
	mem[2421] = 4'b1100;
	mem[2422] = 4'b1100;
	mem[2423] = 4'b1100;
	mem[2424] = 4'b1100;
	mem[2425] = 4'b1100;
	mem[2426] = 4'b0010;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0000;
	mem[2436] = 4'b0000;
	mem[2437] = 4'b0000;
	mem[2438] = 4'b0000;
	mem[2439] = 4'b0000;
	mem[2440] = 4'b0000;
	mem[2441] = 4'b0000;
	mem[2442] = 4'b0000;
	mem[2443] = 4'b0000;
	mem[2444] = 4'b0000;
	mem[2445] = 4'b0000;
	mem[2446] = 4'b0000;
	mem[2447] = 4'b0000;
	mem[2448] = 4'b0000;
	mem[2449] = 4'b0000;
	mem[2450] = 4'b0000;
	mem[2451] = 4'b0000;
	mem[2452] = 4'b0000;
	mem[2453] = 4'b0000;
	mem[2454] = 4'b0000;
	mem[2455] = 4'b0000;
	mem[2456] = 4'b0000;
	mem[2457] = 4'b0000;
	mem[2458] = 4'b0000;
	mem[2459] = 4'b0000;
	mem[2460] = 4'b0000;
	mem[2461] = 4'b0000;
	mem[2462] = 4'b0000;
	mem[2463] = 4'b0000;
	mem[2464] = 4'b0000;
	mem[2465] = 4'b0000;
	mem[2466] = 4'b0000;
	mem[2467] = 4'b0000;
	mem[2468] = 4'b0000;
	mem[2469] = 4'b1010;
	mem[2470] = 4'b1101;
	mem[2471] = 4'b1101;
	mem[2472] = 4'b1101;
	mem[2473] = 4'b1111;
	mem[2474] = 4'b1111;
	mem[2475] = 4'b1111;
	mem[2476] = 4'b1111;
	mem[2477] = 4'b1111;
	mem[2478] = 4'b1111;
	mem[2479] = 4'b1111;
	mem[2480] = 4'b1111;
	mem[2481] = 4'b1101;
	mem[2482] = 4'b1101;
	mem[2483] = 4'b1101;
	mem[2484] = 4'b1101;
	mem[2485] = 4'b1101;
	mem[2486] = 4'b0110;
	mem[2487] = 4'b0000;
	mem[2488] = 4'b0000;
	mem[2489] = 4'b0000;
	mem[2490] = 4'b0000;
	mem[2491] = 4'b0000;
	mem[2492] = 4'b0000;
	mem[2493] = 4'b0000;
	mem[2494] = 4'b0000;
	mem[2495] = 4'b0000;
	mem[2496] = 4'b0000;
	mem[2497] = 4'b0000;
	mem[2498] = 4'b0000;
	mem[2499] = 4'b0000;
	mem[2500] = 4'b0000;
	mem[2501] = 4'b0000;
	mem[2502] = 4'b0000;
	mem[2503] = 4'b0000;
	mem[2504] = 4'b0000;
	mem[2505] = 4'b0000;
	mem[2506] = 4'b0000;
	mem[2507] = 4'b0000;
	mem[2508] = 4'b0000;
	mem[2509] = 4'b0000;
	mem[2510] = 4'b0000;
	mem[2511] = 4'b0000;
	mem[2512] = 4'b0000;
	mem[2513] = 4'b0000;
	mem[2514] = 4'b0000;
	mem[2515] = 4'b0000;
	mem[2516] = 4'b0000;
	mem[2517] = 4'b0000;
	mem[2518] = 4'b0000;
	mem[2519] = 4'b0000;
	mem[2520] = 4'b0000;
	mem[2521] = 4'b0000;
	mem[2522] = 4'b0000;
	mem[2523] = 4'b0000;
	mem[2524] = 4'b0000;
	mem[2525] = 4'b0000;
	mem[2526] = 4'b0000;
	mem[2527] = 4'b0000;
	mem[2528] = 4'b0000;
	mem[2529] = 4'b0000;
	mem[2530] = 4'b0000;
	mem[2531] = 4'b0000;
	mem[2532] = 4'b0001;
	mem[2533] = 4'b0001;
	mem[2534] = 4'b0000;
	mem[2535] = 4'b0000;
	mem[2536] = 4'b0000;
	mem[2537] = 4'b1000;
	mem[2538] = 4'b1100;
	mem[2539] = 4'b1100;
	mem[2540] = 4'b1100;
	mem[2541] = 4'b1100;
	mem[2542] = 4'b1100;
	mem[2543] = 4'b1100;
	mem[2544] = 4'b1100;
	mem[2545] = 4'b1100;
	mem[2546] = 4'b1100;
	mem[2547] = 4'b1100;
	mem[2548] = 4'b1100;
	mem[2549] = 4'b1100;
	mem[2550] = 4'b1100;
	mem[2551] = 4'b1100;
	mem[2552] = 4'b1100;
	mem[2553] = 4'b1100;
	mem[2554] = 4'b0010;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b1000;
	mem[2564] = 4'b1101;
	mem[2565] = 4'b1101;
	mem[2566] = 4'b1101;
	mem[2567] = 4'b1101;
	mem[2568] = 4'b1101;
	mem[2569] = 4'b1100;
	mem[2570] = 4'b1100;
	mem[2571] = 4'b1100;
	mem[2572] = 4'b1100;
	mem[2573] = 4'b1100;
	mem[2574] = 4'b1011;
	mem[2575] = 4'b1011;
	mem[2576] = 4'b1011;
	mem[2577] = 4'b1011;
	mem[2578] = 4'b1011;
	mem[2579] = 4'b1010;
	mem[2580] = 4'b1010;
	mem[2581] = 4'b1010;
	mem[2582] = 4'b1010;
	mem[2583] = 4'b1010;
	mem[2584] = 4'b1001;
	mem[2585] = 4'b1001;
	mem[2586] = 4'b1001;
	mem[2587] = 4'b1001;
	mem[2588] = 4'b1001;
	mem[2589] = 4'b1000;
	mem[2590] = 4'b1000;
	mem[2591] = 4'b1000;
	mem[2592] = 4'b1000;
	mem[2593] = 4'b1000;
	mem[2594] = 4'b0111;
	mem[2595] = 4'b1000;
	mem[2596] = 4'b0111;
	mem[2597] = 4'b0111;
	mem[2598] = 4'b1000;
	mem[2599] = 4'b1000;
	mem[2600] = 4'b0111;
	mem[2601] = 4'b1000;
	mem[2602] = 4'b1000;
	mem[2603] = 4'b1000;
	mem[2604] = 4'b1000;
	mem[2605] = 4'b0111;
	mem[2606] = 4'b0111;
	mem[2607] = 4'b0111;
	mem[2608] = 4'b0111;
	mem[2609] = 4'b0111;
	mem[2610] = 4'b0110;
	mem[2611] = 4'b0110;
	mem[2612] = 4'b0101;
	mem[2613] = 4'b0101;
	mem[2614] = 4'b0100;
	mem[2615] = 4'b0100;
	mem[2616] = 4'b0011;
	mem[2617] = 4'b0011;
	mem[2618] = 4'b0011;
	mem[2619] = 4'b0011;
	mem[2620] = 4'b0010;
	mem[2621] = 4'b0010;
	mem[2622] = 4'b0010;
	mem[2623] = 4'b0010;
	mem[2624] = 4'b0010;
	mem[2625] = 4'b0001;
	mem[2626] = 4'b0001;
	mem[2627] = 4'b0001;
	mem[2628] = 4'b0001;
	mem[2629] = 4'b0001;
	mem[2630] = 4'b0001;
	mem[2631] = 4'b0000;
	mem[2632] = 4'b0000;
	mem[2633] = 4'b0000;
	mem[2634] = 4'b0000;
	mem[2635] = 4'b1000;
	mem[2636] = 4'b1101;
	mem[2637] = 4'b1101;
	mem[2638] = 4'b1101;
	mem[2639] = 4'b1100;
	mem[2640] = 4'b1100;
	mem[2641] = 4'b1100;
	mem[2642] = 4'b1011;
	mem[2643] = 4'b1011;
	mem[2644] = 4'b1011;
	mem[2645] = 4'b1010;
	mem[2646] = 4'b1010;
	mem[2647] = 4'b1010;
	mem[2648] = 4'b1010;
	mem[2649] = 4'b1001;
	mem[2650] = 4'b1001;
	mem[2651] = 4'b1001;
	mem[2652] = 4'b1001;
	mem[2653] = 4'b1000;
	mem[2654] = 4'b0111;
	mem[2655] = 4'b0111;
	mem[2656] = 4'b0111;
	mem[2657] = 4'b0110;
	mem[2658] = 4'b0110;
	mem[2659] = 4'b0111;
	mem[2660] = 4'b0111;
	mem[2661] = 4'b0110;
	mem[2662] = 4'b0101;
	mem[2663] = 4'b0101;
	mem[2664] = 4'b0101;
	mem[2665] = 4'b0110;
	mem[2666] = 4'b0110;
	mem[2667] = 4'b0110;
	mem[2668] = 4'b0101;
	mem[2669] = 4'b0101;
	mem[2670] = 4'b0101;
	mem[2671] = 4'b0101;
	mem[2672] = 4'b0100;
	mem[2673] = 4'b0100;
	mem[2674] = 4'b0100;
	mem[2675] = 4'b0100;
	mem[2676] = 4'b0011;
	mem[2677] = 4'b0011;
	mem[2678] = 4'b0011;
	mem[2679] = 4'b0011;
	mem[2680] = 4'b0011;
	mem[2681] = 4'b0010;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b1001;
	mem[2692] = 4'b1111;
	mem[2693] = 4'b1111;
	mem[2694] = 4'b1111;
	mem[2695] = 4'b1111;
	mem[2696] = 4'b1110;
	mem[2697] = 4'b1110;
	mem[2698] = 4'b1110;
	mem[2699] = 4'b1110;
	mem[2700] = 4'b1101;
	mem[2701] = 4'b1101;
	mem[2702] = 4'b1101;
	mem[2703] = 4'b1101;
	mem[2704] = 4'b1101;
	mem[2705] = 4'b1100;
	mem[2706] = 4'b1100;
	mem[2707] = 4'b1100;
	mem[2708] = 4'b1100;
	mem[2709] = 4'b1011;
	mem[2710] = 4'b1011;
	mem[2711] = 4'b1011;
	mem[2712] = 4'b1011;
	mem[2713] = 4'b1011;
	mem[2714] = 4'b1010;
	mem[2715] = 4'b1010;
	mem[2716] = 4'b1010;
	mem[2717] = 4'b1010;
	mem[2718] = 4'b1001;
	mem[2719] = 4'b1001;
	mem[2720] = 4'b1001;
	mem[2721] = 4'b1001;
	mem[2722] = 4'b1001;
	mem[2723] = 4'b1000;
	mem[2724] = 4'b1000;
	mem[2725] = 4'b0111;
	mem[2726] = 4'b0111;
	mem[2727] = 4'b0111;
	mem[2728] = 4'b0111;
	mem[2729] = 4'b0110;
	mem[2730] = 4'b0111;
	mem[2731] = 4'b0111;
	mem[2732] = 4'b0110;
	mem[2733] = 4'b0110;
	mem[2734] = 4'b0110;
	mem[2735] = 4'b0110;
	mem[2736] = 4'b0101;
	mem[2737] = 4'b0101;
	mem[2738] = 4'b0101;
	mem[2739] = 4'b0100;
	mem[2740] = 4'b0100;
	mem[2741] = 4'b0100;
	mem[2742] = 4'b0100;
	mem[2743] = 4'b0101;
	mem[2744] = 4'b0100;
	mem[2745] = 4'b0100;
	mem[2746] = 4'b0011;
	mem[2747] = 4'b0011;
	mem[2748] = 4'b0011;
	mem[2749] = 4'b0011;
	mem[2750] = 4'b0010;
	mem[2751] = 4'b0010;
	mem[2752] = 4'b0010;
	mem[2753] = 4'b0010;
	mem[2754] = 4'b0010;
	mem[2755] = 4'b0001;
	mem[2756] = 4'b0001;
	mem[2757] = 4'b0001;
	mem[2758] = 4'b0001;
	mem[2759] = 4'b0000;
	mem[2760] = 4'b0000;
	mem[2761] = 4'b0000;
	mem[2762] = 4'b0000;
	mem[2763] = 4'b1001;
	mem[2764] = 4'b1111;
	mem[2765] = 4'b1111;
	mem[2766] = 4'b1110;
	mem[2767] = 4'b1110;
	mem[2768] = 4'b1110;
	mem[2769] = 4'b1101;
	mem[2770] = 4'b1101;
	mem[2771] = 4'b1101;
	mem[2772] = 4'b1100;
	mem[2773] = 4'b1100;
	mem[2774] = 4'b1100;
	mem[2775] = 4'b1011;
	mem[2776] = 4'b1011;
	mem[2777] = 4'b1011;
	mem[2778] = 4'b1010;
	mem[2779] = 4'b1001;
	mem[2780] = 4'b1010;
	mem[2781] = 4'b1001;
	mem[2782] = 4'b1001;
	mem[2783] = 4'b1000;
	mem[2784] = 4'b0111;
	mem[2785] = 4'b0111;
	mem[2786] = 4'b1000;
	mem[2787] = 4'b1000;
	mem[2788] = 4'b0111;
	mem[2789] = 4'b0111;
	mem[2790] = 4'b0110;
	mem[2791] = 4'b0110;
	mem[2792] = 4'b0110;
	mem[2793] = 4'b0101;
	mem[2794] = 4'b0101;
	mem[2795] = 4'b0101;
	mem[2796] = 4'b0100;
	mem[2797] = 4'b0100;
	mem[2798] = 4'b0100;
	mem[2799] = 4'b0100;
	mem[2800] = 4'b0011;
	mem[2801] = 4'b0011;
	mem[2802] = 4'b0011;
	mem[2803] = 4'b0011;
	mem[2804] = 4'b0010;
	mem[2805] = 4'b0010;
	mem[2806] = 4'b0010;
	mem[2807] = 4'b0010;
	mem[2808] = 4'b0010;
	mem[2809] = 4'b0001;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b1001;
	mem[2820] = 4'b1111;
	mem[2821] = 4'b1111;
	mem[2822] = 4'b1111;
	mem[2823] = 4'b1111;
	mem[2824] = 4'b1110;
	mem[2825] = 4'b1110;
	mem[2826] = 4'b1110;
	mem[2827] = 4'b1110;
	mem[2828] = 4'b1101;
	mem[2829] = 4'b1101;
	mem[2830] = 4'b1101;
	mem[2831] = 4'b1101;
	mem[2832] = 4'b1101;
	mem[2833] = 4'b1100;
	mem[2834] = 4'b1100;
	mem[2835] = 4'b1100;
	mem[2836] = 4'b1100;
	mem[2837] = 4'b1011;
	mem[2838] = 4'b1011;
	mem[2839] = 4'b1011;
	mem[2840] = 4'b1011;
	mem[2841] = 4'b1011;
	mem[2842] = 4'b1010;
	mem[2843] = 4'b1010;
	mem[2844] = 4'b1010;
	mem[2845] = 4'b1010;
	mem[2846] = 4'b1001;
	mem[2847] = 4'b1001;
	mem[2848] = 4'b1001;
	mem[2849] = 4'b1001;
	mem[2850] = 4'b1001;
	mem[2851] = 4'b1000;
	mem[2852] = 4'b1000;
	mem[2853] = 4'b1000;
	mem[2854] = 4'b0111;
	mem[2855] = 4'b0111;
	mem[2856] = 4'b0111;
	mem[2857] = 4'b0110;
	mem[2858] = 4'b0110;
	mem[2859] = 4'b0111;
	mem[2860] = 4'b0111;
	mem[2861] = 4'b0110;
	mem[2862] = 4'b0110;
	mem[2863] = 4'b0110;
	mem[2864] = 4'b0101;
	mem[2865] = 4'b0101;
	mem[2866] = 4'b0101;
	mem[2867] = 4'b0101;
	mem[2868] = 4'b0100;
	mem[2869] = 4'b0100;
	mem[2870] = 4'b0101;
	mem[2871] = 4'b0100;
	mem[2872] = 4'b0100;
	mem[2873] = 4'b0100;
	mem[2874] = 4'b0011;
	mem[2875] = 4'b0011;
	mem[2876] = 4'b0011;
	mem[2877] = 4'b0011;
	mem[2878] = 4'b0010;
	mem[2879] = 4'b0010;
	mem[2880] = 4'b0010;
	mem[2881] = 4'b0010;
	mem[2882] = 4'b0010;
	mem[2883] = 4'b0001;
	mem[2884] = 4'b0001;
	mem[2885] = 4'b0001;
	mem[2886] = 4'b0001;
	mem[2887] = 4'b0000;
	mem[2888] = 4'b0000;
	mem[2889] = 4'b0000;
	mem[2890] = 4'b0000;
	mem[2891] = 4'b1001;
	mem[2892] = 4'b1111;
	mem[2893] = 4'b1111;
	mem[2894] = 4'b1110;
	mem[2895] = 4'b1110;
	mem[2896] = 4'b1110;
	mem[2897] = 4'b1101;
	mem[2898] = 4'b1101;
	mem[2899] = 4'b1101;
	mem[2900] = 4'b1100;
	mem[2901] = 4'b1100;
	mem[2902] = 4'b1100;
	mem[2903] = 4'b1011;
	mem[2904] = 4'b1011;
	mem[2905] = 4'b1010;
	mem[2906] = 4'b1001;
	mem[2907] = 4'b1001;
	mem[2908] = 4'b1001;
	mem[2909] = 4'b1010;
	mem[2910] = 4'b1001;
	mem[2911] = 4'b1000;
	mem[2912] = 4'b0111;
	mem[2913] = 4'b1000;
	mem[2914] = 4'b1000;
	mem[2915] = 4'b0111;
	mem[2916] = 4'b0111;
	mem[2917] = 4'b0111;
	mem[2918] = 4'b0110;
	mem[2919] = 4'b0110;
	mem[2920] = 4'b0110;
	mem[2921] = 4'b0101;
	mem[2922] = 4'b0101;
	mem[2923] = 4'b0101;
	mem[2924] = 4'b0101;
	mem[2925] = 4'b0100;
	mem[2926] = 4'b0100;
	mem[2927] = 4'b0100;
	mem[2928] = 4'b0100;
	mem[2929] = 4'b0011;
	mem[2930] = 4'b0011;
	mem[2931] = 4'b0011;
	mem[2932] = 4'b0011;
	mem[2933] = 4'b0010;
	mem[2934] = 4'b0010;
	mem[2935] = 4'b0010;
	mem[2936] = 4'b0010;
	mem[2937] = 4'b0010;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b1001;
	mem[2948] = 4'b1111;
	mem[2949] = 4'b1111;
	mem[2950] = 4'b1111;
	mem[2951] = 4'b1111;
	mem[2952] = 4'b1110;
	mem[2953] = 4'b1110;
	mem[2954] = 4'b1110;
	mem[2955] = 4'b1110;
	mem[2956] = 4'b1101;
	mem[2957] = 4'b1101;
	mem[2958] = 4'b1101;
	mem[2959] = 4'b1101;
	mem[2960] = 4'b1101;
	mem[2961] = 4'b1100;
	mem[2962] = 4'b1100;
	mem[2963] = 4'b1100;
	mem[2964] = 4'b1100;
	mem[2965] = 4'b1011;
	mem[2966] = 4'b1011;
	mem[2967] = 4'b1011;
	mem[2968] = 4'b1011;
	mem[2969] = 4'b1011;
	mem[2970] = 4'b1010;
	mem[2971] = 4'b1010;
	mem[2972] = 4'b1010;
	mem[2973] = 4'b1010;
	mem[2974] = 4'b1001;
	mem[2975] = 4'b1001;
	mem[2976] = 4'b1001;
	mem[2977] = 4'b1001;
	mem[2978] = 4'b1001;
	mem[2979] = 4'b1000;
	mem[2980] = 4'b1000;
	mem[2981] = 4'b1000;
	mem[2982] = 4'b1000;
	mem[2983] = 4'b0111;
	mem[2984] = 4'b0110;
	mem[2985] = 4'b0110;
	mem[2986] = 4'b0110;
	mem[2987] = 4'b0110;
	mem[2988] = 4'b0111;
	mem[2989] = 4'b0110;
	mem[2990] = 4'b0110;
	mem[2991] = 4'b0110;
	mem[2992] = 4'b0101;
	mem[2993] = 4'b0101;
	mem[2994] = 4'b0101;
	mem[2995] = 4'b0101;
	mem[2996] = 4'b0101;
	mem[2997] = 4'b0101;
	mem[2998] = 4'b0101;
	mem[2999] = 4'b0100;
	mem[3000] = 4'b0100;
	mem[3001] = 4'b0100;
	mem[3002] = 4'b0011;
	mem[3003] = 4'b0011;
	mem[3004] = 4'b0011;
	mem[3005] = 4'b0011;
	mem[3006] = 4'b0010;
	mem[3007] = 4'b0010;
	mem[3008] = 4'b0010;
	mem[3009] = 4'b0010;
	mem[3010] = 4'b0010;
	mem[3011] = 4'b0001;
	mem[3012] = 4'b0001;
	mem[3013] = 4'b0001;
	mem[3014] = 4'b0001;
	mem[3015] = 4'b0000;
	mem[3016] = 4'b0000;
	mem[3017] = 4'b0000;
	mem[3018] = 4'b0000;
	mem[3019] = 4'b1001;
	mem[3020] = 4'b1111;
	mem[3021] = 4'b1111;
	mem[3022] = 4'b1110;
	mem[3023] = 4'b1110;
	mem[3024] = 4'b1110;
	mem[3025] = 4'b1101;
	mem[3026] = 4'b1101;
	mem[3027] = 4'b1101;
	mem[3028] = 4'b1100;
	mem[3029] = 4'b1100;
	mem[3030] = 4'b1100;
	mem[3031] = 4'b1011;
	mem[3032] = 4'b1010;
	mem[3033] = 4'b1001;
	mem[3034] = 4'b1001;
	mem[3035] = 4'b1001;
	mem[3036] = 4'b1010;
	mem[3037] = 4'b1010;
	mem[3038] = 4'b1001;
	mem[3039] = 4'b1001;
	mem[3040] = 4'b1001;
	mem[3041] = 4'b1001;
	mem[3042] = 4'b1000;
	mem[3043] = 4'b0111;
	mem[3044] = 4'b0111;
	mem[3045] = 4'b0111;
	mem[3046] = 4'b0110;
	mem[3047] = 4'b0110;
	mem[3048] = 4'b0110;
	mem[3049] = 4'b0110;
	mem[3050] = 4'b0101;
	mem[3051] = 4'b0101;
	mem[3052] = 4'b0101;
	mem[3053] = 4'b0101;
	mem[3054] = 4'b0100;
	mem[3055] = 4'b0100;
	mem[3056] = 4'b0100;
	mem[3057] = 4'b0100;
	mem[3058] = 4'b0011;
	mem[3059] = 4'b0011;
	mem[3060] = 4'b0011;
	mem[3061] = 4'b0011;
	mem[3062] = 4'b0011;
	mem[3063] = 4'b0010;
	mem[3064] = 4'b0010;
	mem[3065] = 4'b0010;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b1001;
	mem[3076] = 4'b1111;
	mem[3077] = 4'b1111;
	mem[3078] = 4'b1111;
	mem[3079] = 4'b1111;
	mem[3080] = 4'b1110;
	mem[3081] = 4'b1110;
	mem[3082] = 4'b1110;
	mem[3083] = 4'b1110;
	mem[3084] = 4'b1101;
	mem[3085] = 4'b1101;
	mem[3086] = 4'b1101;
	mem[3087] = 4'b1101;
	mem[3088] = 4'b1101;
	mem[3089] = 4'b1100;
	mem[3090] = 4'b1100;
	mem[3091] = 4'b1100;
	mem[3092] = 4'b1100;
	mem[3093] = 4'b1011;
	mem[3094] = 4'b1011;
	mem[3095] = 4'b1011;
	mem[3096] = 4'b1011;
	mem[3097] = 4'b1011;
	mem[3098] = 4'b1010;
	mem[3099] = 4'b1010;
	mem[3100] = 4'b1010;
	mem[3101] = 4'b1010;
	mem[3102] = 4'b1001;
	mem[3103] = 4'b1001;
	mem[3104] = 4'b1001;
	mem[3105] = 4'b1001;
	mem[3106] = 4'b1001;
	mem[3107] = 4'b1000;
	mem[3108] = 4'b1000;
	mem[3109] = 4'b1000;
	mem[3110] = 4'b1000;
	mem[3111] = 4'b1000;
	mem[3112] = 4'b0111;
	mem[3113] = 4'b0110;
	mem[3114] = 4'b0110;
	mem[3115] = 4'b0110;
	mem[3116] = 4'b0110;
	mem[3117] = 4'b0110;
	mem[3118] = 4'b0110;
	mem[3119] = 4'b0110;
	mem[3120] = 4'b0101;
	mem[3121] = 4'b0101;
	mem[3122] = 4'b0101;
	mem[3123] = 4'b0101;
	mem[3124] = 4'b0101;
	mem[3125] = 4'b0101;
	mem[3126] = 4'b0100;
	mem[3127] = 4'b0100;
	mem[3128] = 4'b0100;
	mem[3129] = 4'b0100;
	mem[3130] = 4'b0011;
	mem[3131] = 4'b0011;
	mem[3132] = 4'b0011;
	mem[3133] = 4'b0011;
	mem[3134] = 4'b0010;
	mem[3135] = 4'b0010;
	mem[3136] = 4'b0010;
	mem[3137] = 4'b0010;
	mem[3138] = 4'b0010;
	mem[3139] = 4'b0001;
	mem[3140] = 4'b0001;
	mem[3141] = 4'b0001;
	mem[3142] = 4'b0001;
	mem[3143] = 4'b0000;
	mem[3144] = 4'b0000;
	mem[3145] = 4'b0000;
	mem[3146] = 4'b0000;
	mem[3147] = 4'b1001;
	mem[3148] = 4'b1111;
	mem[3149] = 4'b1111;
	mem[3150] = 4'b1110;
	mem[3151] = 4'b1110;
	mem[3152] = 4'b1110;
	mem[3153] = 4'b1101;
	mem[3154] = 4'b1101;
	mem[3155] = 4'b1100;
	mem[3156] = 4'b1011;
	mem[3157] = 4'b1011;
	mem[3158] = 4'b1100;
	mem[3159] = 4'b1011;
	mem[3160] = 4'b1011;
	mem[3161] = 4'b1001;
	mem[3162] = 4'b1001;
	mem[3163] = 4'b1011;
	mem[3164] = 4'b1010;
	mem[3165] = 4'b1001;
	mem[3166] = 4'b1001;
	mem[3167] = 4'b1001;
	mem[3168] = 4'b1000;
	mem[3169] = 4'b1000;
	mem[3170] = 4'b1000;
	mem[3171] = 4'b0111;
	mem[3172] = 4'b0111;
	mem[3173] = 4'b0111;
	mem[3174] = 4'b0110;
	mem[3175] = 4'b0110;
	mem[3176] = 4'b0110;
	mem[3177] = 4'b0110;
	mem[3178] = 4'b0101;
	mem[3179] = 4'b0101;
	mem[3180] = 4'b0101;
	mem[3181] = 4'b0101;
	mem[3182] = 4'b0100;
	mem[3183] = 4'b0100;
	mem[3184] = 4'b0100;
	mem[3185] = 4'b0100;
	mem[3186] = 4'b0100;
	mem[3187] = 4'b0011;
	mem[3188] = 4'b0011;
	mem[3189] = 4'b0011;
	mem[3190] = 4'b0011;
	mem[3191] = 4'b0011;
	mem[3192] = 4'b0010;
	mem[3193] = 4'b0010;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b1001;
	mem[3204] = 4'b1111;
	mem[3205] = 4'b1111;
	mem[3206] = 4'b1111;
	mem[3207] = 4'b1111;
	mem[3208] = 4'b1110;
	mem[3209] = 4'b1110;
	mem[3210] = 4'b1110;
	mem[3211] = 4'b1110;
	mem[3212] = 4'b1101;
	mem[3213] = 4'b1101;
	mem[3214] = 4'b1101;
	mem[3215] = 4'b1101;
	mem[3216] = 4'b1101;
	mem[3217] = 4'b1100;
	mem[3218] = 4'b1100;
	mem[3219] = 4'b1100;
	mem[3220] = 4'b1100;
	mem[3221] = 4'b1011;
	mem[3222] = 4'b1011;
	mem[3223] = 4'b1011;
	mem[3224] = 4'b1011;
	mem[3225] = 4'b1011;
	mem[3226] = 4'b1010;
	mem[3227] = 4'b1010;
	mem[3228] = 4'b1010;
	mem[3229] = 4'b1001;
	mem[3230] = 4'b1001;
	mem[3231] = 4'b1000;
	mem[3232] = 4'b1000;
	mem[3233] = 4'b1000;
	mem[3234] = 4'b1000;
	mem[3235] = 4'b1000;
	mem[3236] = 4'b1000;
	mem[3237] = 4'b1000;
	mem[3238] = 4'b1000;
	mem[3239] = 4'b0111;
	mem[3240] = 4'b1000;
	mem[3241] = 4'b0110;
	mem[3242] = 4'b0110;
	mem[3243] = 4'b0110;
	mem[3244] = 4'b0110;
	mem[3245] = 4'b0101;
	mem[3246] = 4'b0110;
	mem[3247] = 4'b0110;
	mem[3248] = 4'b0101;
	mem[3249] = 4'b0101;
	mem[3250] = 4'b0101;
	mem[3251] = 4'b0101;
	mem[3252] = 4'b0101;
	mem[3253] = 4'b0100;
	mem[3254] = 4'b0100;
	mem[3255] = 4'b0100;
	mem[3256] = 4'b0100;
	mem[3257] = 4'b0100;
	mem[3258] = 4'b0011;
	mem[3259] = 4'b0011;
	mem[3260] = 4'b0011;
	mem[3261] = 4'b0011;
	mem[3262] = 4'b0010;
	mem[3263] = 4'b0010;
	mem[3264] = 4'b0010;
	mem[3265] = 4'b0010;
	mem[3266] = 4'b0010;
	mem[3267] = 4'b0001;
	mem[3268] = 4'b0001;
	mem[3269] = 4'b0001;
	mem[3270] = 4'b0001;
	mem[3271] = 4'b0000;
	mem[3272] = 4'b0000;
	mem[3273] = 4'b0000;
	mem[3274] = 4'b0000;
	mem[3275] = 4'b1001;
	mem[3276] = 4'b1111;
	mem[3277] = 4'b1111;
	mem[3278] = 4'b1110;
	mem[3279] = 4'b1110;
	mem[3280] = 4'b1110;
	mem[3281] = 4'b1101;
	mem[3282] = 4'b1100;
	mem[3283] = 4'b1011;
	mem[3284] = 4'b1011;
	mem[3285] = 4'b1100;
	mem[3286] = 4'b1100;
	mem[3287] = 4'b1011;
	mem[3288] = 4'b1011;
	mem[3289] = 4'b1011;
	mem[3290] = 4'b1011;
	mem[3291] = 4'b1010;
	mem[3292] = 4'b1010;
	mem[3293] = 4'b1001;
	mem[3294] = 4'b1001;
	mem[3295] = 4'b1001;
	mem[3296] = 4'b1000;
	mem[3297] = 4'b1000;
	mem[3298] = 4'b1000;
	mem[3299] = 4'b0111;
	mem[3300] = 4'b0111;
	mem[3301] = 4'b0111;
	mem[3302] = 4'b0111;
	mem[3303] = 4'b0110;
	mem[3304] = 4'b0110;
	mem[3305] = 4'b0110;
	mem[3306] = 4'b0110;
	mem[3307] = 4'b0101;
	mem[3308] = 4'b0101;
	mem[3309] = 4'b0101;
	mem[3310] = 4'b0101;
	mem[3311] = 4'b0100;
	mem[3312] = 4'b0100;
	mem[3313] = 4'b0100;
	mem[3314] = 4'b0100;
	mem[3315] = 4'b0100;
	mem[3316] = 4'b0011;
	mem[3317] = 4'b0011;
	mem[3318] = 4'b0011;
	mem[3319] = 4'b0011;
	mem[3320] = 4'b0011;
	mem[3321] = 4'b0010;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b1001;
	mem[3332] = 4'b1111;
	mem[3333] = 4'b1111;
	mem[3334] = 4'b1111;
	mem[3335] = 4'b1111;
	mem[3336] = 4'b1110;
	mem[3337] = 4'b1110;
	mem[3338] = 4'b1110;
	mem[3339] = 4'b1110;
	mem[3340] = 4'b1101;
	mem[3341] = 4'b1101;
	mem[3342] = 4'b1101;
	mem[3343] = 4'b1101;
	mem[3344] = 4'b1101;
	mem[3345] = 4'b1100;
	mem[3346] = 4'b1100;
	mem[3347] = 4'b1100;
	mem[3348] = 4'b1100;
	mem[3349] = 4'b1011;
	mem[3350] = 4'b1011;
	mem[3351] = 4'b1011;
	mem[3352] = 4'b1011;
	mem[3353] = 4'b1011;
	mem[3354] = 4'b1010;
	mem[3355] = 4'b1010;
	mem[3356] = 4'b1001;
	mem[3357] = 4'b1001;
	mem[3358] = 4'b1000;
	mem[3359] = 4'b1000;
	mem[3360] = 4'b1000;
	mem[3361] = 4'b1000;
	mem[3362] = 4'b1000;
	mem[3363] = 4'b0111;
	mem[3364] = 4'b0111;
	mem[3365] = 4'b1000;
	mem[3366] = 4'b1000;
	mem[3367] = 4'b0111;
	mem[3368] = 4'b0111;
	mem[3369] = 4'b0111;
	mem[3370] = 4'b0110;
	mem[3371] = 4'b0110;
	mem[3372] = 4'b0110;
	mem[3373] = 4'b0110;
	mem[3374] = 4'b0101;
	mem[3375] = 4'b0110;
	mem[3376] = 4'b0110;
	mem[3377] = 4'b0101;
	mem[3378] = 4'b0101;
	mem[3379] = 4'b0101;
	mem[3380] = 4'b0101;
	mem[3381] = 4'b0100;
	mem[3382] = 4'b0100;
	mem[3383] = 4'b0100;
	mem[3384] = 4'b0100;
	mem[3385] = 4'b0100;
	mem[3386] = 4'b0011;
	mem[3387] = 4'b0011;
	mem[3388] = 4'b0011;
	mem[3389] = 4'b0011;
	mem[3390] = 4'b0010;
	mem[3391] = 4'b0010;
	mem[3392] = 4'b0010;
	mem[3393] = 4'b0010;
	mem[3394] = 4'b0010;
	mem[3395] = 4'b0001;
	mem[3396] = 4'b0001;
	mem[3397] = 4'b0001;
	mem[3398] = 4'b0001;
	mem[3399] = 4'b0000;
	mem[3400] = 4'b0000;
	mem[3401] = 4'b0000;
	mem[3402] = 4'b0000;
	mem[3403] = 4'b1001;
	mem[3404] = 4'b1111;
	mem[3405] = 4'b1111;
	mem[3406] = 4'b1110;
	mem[3407] = 4'b1110;
	mem[3408] = 4'b1110;
	mem[3409] = 4'b1100;
	mem[3410] = 4'b1011;
	mem[3411] = 4'b1100;
	mem[3412] = 4'b1100;
	mem[3413] = 4'b1100;
	mem[3414] = 4'b1011;
	mem[3415] = 4'b1010;
	mem[3416] = 4'b1011;
	mem[3417] = 4'b1011;
	mem[3418] = 4'b1010;
	mem[3419] = 4'b1010;
	mem[3420] = 4'b1010;
	mem[3421] = 4'b1001;
	mem[3422] = 4'b1001;
	mem[3423] = 4'b1001;
	mem[3424] = 4'b1000;
	mem[3425] = 4'b1000;
	mem[3426] = 4'b1000;
	mem[3427] = 4'b1000;
	mem[3428] = 4'b0111;
	mem[3429] = 4'b0111;
	mem[3430] = 4'b0111;
	mem[3431] = 4'b0111;
	mem[3432] = 4'b0110;
	mem[3433] = 4'b0110;
	mem[3434] = 4'b0110;
	mem[3435] = 4'b0110;
	mem[3436] = 4'b0101;
	mem[3437] = 4'b0101;
	mem[3438] = 4'b0101;
	mem[3439] = 4'b0101;
	mem[3440] = 4'b0100;
	mem[3441] = 4'b0100;
	mem[3442] = 4'b0100;
	mem[3443] = 4'b0100;
	mem[3444] = 4'b0100;
	mem[3445] = 4'b0011;
	mem[3446] = 4'b0011;
	mem[3447] = 4'b0011;
	mem[3448] = 4'b0011;
	mem[3449] = 4'b0011;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b1001;
	mem[3460] = 4'b1111;
	mem[3461] = 4'b1111;
	mem[3462] = 4'b1111;
	mem[3463] = 4'b1111;
	mem[3464] = 4'b1110;
	mem[3465] = 4'b1110;
	mem[3466] = 4'b1110;
	mem[3467] = 4'b1110;
	mem[3468] = 4'b1101;
	mem[3469] = 4'b1101;
	mem[3470] = 4'b1101;
	mem[3471] = 4'b1101;
	mem[3472] = 4'b1101;
	mem[3473] = 4'b1100;
	mem[3474] = 4'b1100;
	mem[3475] = 4'b1100;
	mem[3476] = 4'b1100;
	mem[3477] = 4'b1011;
	mem[3478] = 4'b1011;
	mem[3479] = 4'b1011;
	mem[3480] = 4'b1011;
	mem[3481] = 4'b1011;
	mem[3482] = 4'b1010;
	mem[3483] = 4'b1001;
	mem[3484] = 4'b1001;
	mem[3485] = 4'b1001;
	mem[3486] = 4'b1000;
	mem[3487] = 4'b1000;
	mem[3488] = 4'b1000;
	mem[3489] = 4'b1000;
	mem[3490] = 4'b1000;
	mem[3491] = 4'b0111;
	mem[3492] = 4'b0111;
	mem[3493] = 4'b0111;
	mem[3494] = 4'b1000;
	mem[3495] = 4'b1000;
	mem[3496] = 4'b0111;
	mem[3497] = 4'b0111;
	mem[3498] = 4'b0111;
	mem[3499] = 4'b0110;
	mem[3500] = 4'b0110;
	mem[3501] = 4'b0110;
	mem[3502] = 4'b0101;
	mem[3503] = 4'b0101;
	mem[3504] = 4'b0110;
	mem[3505] = 4'b0101;
	mem[3506] = 4'b0101;
	mem[3507] = 4'b0101;
	mem[3508] = 4'b0101;
	mem[3509] = 4'b0100;
	mem[3510] = 4'b0100;
	mem[3511] = 4'b0100;
	mem[3512] = 4'b0100;
	mem[3513] = 4'b0100;
	mem[3514] = 4'b0011;
	mem[3515] = 4'b0011;
	mem[3516] = 4'b0011;
	mem[3517] = 4'b0011;
	mem[3518] = 4'b0010;
	mem[3519] = 4'b0010;
	mem[3520] = 4'b0010;
	mem[3521] = 4'b0010;
	mem[3522] = 4'b0010;
	mem[3523] = 4'b0001;
	mem[3524] = 4'b0001;
	mem[3525] = 4'b0001;
	mem[3526] = 4'b0001;
	mem[3527] = 4'b0000;
	mem[3528] = 4'b0000;
	mem[3529] = 4'b0000;
	mem[3530] = 4'b0000;
	mem[3531] = 4'b1001;
	mem[3532] = 4'b1111;
	mem[3533] = 4'b1111;
	mem[3534] = 4'b1110;
	mem[3535] = 4'b1110;
	mem[3536] = 4'b1101;
	mem[3537] = 4'b1100;
	mem[3538] = 4'b1101;
	mem[3539] = 4'b1101;
	mem[3540] = 4'b1100;
	mem[3541] = 4'b1011;
	mem[3542] = 4'b1010;
	mem[3543] = 4'b1010;
	mem[3544] = 4'b1001;
	mem[3545] = 4'b1011;
	mem[3546] = 4'b1010;
	mem[3547] = 4'b1010;
	mem[3548] = 4'b1010;
	mem[3549] = 4'b1001;
	mem[3550] = 4'b1001;
	mem[3551] = 4'b1001;
	mem[3552] = 4'b1001;
	mem[3553] = 4'b1000;
	mem[3554] = 4'b1000;
	mem[3555] = 4'b1000;
	mem[3556] = 4'b0111;
	mem[3557] = 4'b0111;
	mem[3558] = 4'b0111;
	mem[3559] = 4'b0111;
	mem[3560] = 4'b0110;
	mem[3561] = 4'b0110;
	mem[3562] = 4'b0110;
	mem[3563] = 4'b0110;
	mem[3564] = 4'b0110;
	mem[3565] = 4'b0101;
	mem[3566] = 4'b0101;
	mem[3567] = 4'b0101;
	mem[3568] = 4'b0101;
	mem[3569] = 4'b0100;
	mem[3570] = 4'b0100;
	mem[3571] = 4'b0100;
	mem[3572] = 4'b0100;
	mem[3573] = 4'b0100;
	mem[3574] = 4'b0100;
	mem[3575] = 4'b0011;
	mem[3576] = 4'b0011;
	mem[3577] = 4'b0011;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b1001;
	mem[3588] = 4'b1111;
	mem[3589] = 4'b1111;
	mem[3590] = 4'b1111;
	mem[3591] = 4'b1111;
	mem[3592] = 4'b1110;
	mem[3593] = 4'b1110;
	mem[3594] = 4'b1110;
	mem[3595] = 4'b1110;
	mem[3596] = 4'b1101;
	mem[3597] = 4'b1101;
	mem[3598] = 4'b1101;
	mem[3599] = 4'b1101;
	mem[3600] = 4'b1101;
	mem[3601] = 4'b1100;
	mem[3602] = 4'b1100;
	mem[3603] = 4'b1100;
	mem[3604] = 4'b1100;
	mem[3605] = 4'b1011;
	mem[3606] = 4'b1011;
	mem[3607] = 4'b1011;
	mem[3608] = 4'b1011;
	mem[3609] = 4'b1011;
	mem[3610] = 4'b1010;
	mem[3611] = 4'b1001;
	mem[3612] = 4'b1001;
	mem[3613] = 4'b1001;
	mem[3614] = 4'b1001;
	mem[3615] = 4'b1001;
	mem[3616] = 4'b1001;
	mem[3617] = 4'b1000;
	mem[3618] = 4'b1000;
	mem[3619] = 4'b0111;
	mem[3620] = 4'b0111;
	mem[3621] = 4'b0111;
	mem[3622] = 4'b0111;
	mem[3623] = 4'b1000;
	mem[3624] = 4'b0111;
	mem[3625] = 4'b0111;
	mem[3626] = 4'b0111;
	mem[3627] = 4'b0111;
	mem[3628] = 4'b0110;
	mem[3629] = 4'b0110;
	mem[3630] = 4'b0101;
	mem[3631] = 4'b0101;
	mem[3632] = 4'b0110;
	mem[3633] = 4'b0101;
	mem[3634] = 4'b0101;
	mem[3635] = 4'b0101;
	mem[3636] = 4'b0101;
	mem[3637] = 4'b0100;
	mem[3638] = 4'b0100;
	mem[3639] = 4'b0100;
	mem[3640] = 4'b0100;
	mem[3641] = 4'b0100;
	mem[3642] = 4'b0011;
	mem[3643] = 4'b0011;
	mem[3644] = 4'b0011;
	mem[3645] = 4'b0011;
	mem[3646] = 4'b0010;
	mem[3647] = 4'b0010;
	mem[3648] = 4'b0010;
	mem[3649] = 4'b0010;
	mem[3650] = 4'b0010;
	mem[3651] = 4'b0001;
	mem[3652] = 4'b0001;
	mem[3653] = 4'b0001;
	mem[3654] = 4'b0001;
	mem[3655] = 4'b0000;
	mem[3656] = 4'b0000;
	mem[3657] = 4'b0000;
	mem[3658] = 4'b0000;
	mem[3659] = 4'b1001;
	mem[3660] = 4'b1111;
	mem[3661] = 4'b1111;
	mem[3662] = 4'b1110;
	mem[3663] = 4'b1110;
	mem[3664] = 4'b1101;
	mem[3665] = 4'b1100;
	mem[3666] = 4'b1100;
	mem[3667] = 4'b1100;
	mem[3668] = 4'b1011;
	mem[3669] = 4'b1010;
	mem[3670] = 4'b1010;
	mem[3671] = 4'b1010;
	mem[3672] = 4'b1010;
	mem[3673] = 4'b1010;
	mem[3674] = 4'b1011;
	mem[3675] = 4'b1010;
	mem[3676] = 4'b1010;
	mem[3677] = 4'b1010;
	mem[3678] = 4'b1001;
	mem[3679] = 4'b1001;
	mem[3680] = 4'b1001;
	mem[3681] = 4'b1000;
	mem[3682] = 4'b1000;
	mem[3683] = 4'b1000;
	mem[3684] = 4'b1000;
	mem[3685] = 4'b0111;
	mem[3686] = 4'b0111;
	mem[3687] = 4'b0111;
	mem[3688] = 4'b0111;
	mem[3689] = 4'b0110;
	mem[3690] = 4'b0110;
	mem[3691] = 4'b0110;
	mem[3692] = 4'b0110;
	mem[3693] = 4'b0110;
	mem[3694] = 4'b0101;
	mem[3695] = 4'b0101;
	mem[3696] = 4'b0101;
	mem[3697] = 4'b0101;
	mem[3698] = 4'b0101;
	mem[3699] = 4'b0100;
	mem[3700] = 4'b0100;
	mem[3701] = 4'b0100;
	mem[3702] = 4'b0100;
	mem[3703] = 4'b0100;
	mem[3704] = 4'b0100;
	mem[3705] = 4'b0011;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b1001;
	mem[3716] = 4'b1111;
	mem[3717] = 4'b1111;
	mem[3718] = 4'b1111;
	mem[3719] = 4'b1111;
	mem[3720] = 4'b1110;
	mem[3721] = 4'b1110;
	mem[3722] = 4'b1110;
	mem[3723] = 4'b1110;
	mem[3724] = 4'b1101;
	mem[3725] = 4'b1101;
	mem[3726] = 4'b1101;
	mem[3727] = 4'b1101;
	mem[3728] = 4'b1101;
	mem[3729] = 4'b1100;
	mem[3730] = 4'b1100;
	mem[3731] = 4'b1100;
	mem[3732] = 4'b1100;
	mem[3733] = 4'b1011;
	mem[3734] = 4'b1011;
	mem[3735] = 4'b1011;
	mem[3736] = 4'b1011;
	mem[3737] = 4'b1010;
	mem[3738] = 4'b1001;
	mem[3739] = 4'b1001;
	mem[3740] = 4'b1001;
	mem[3741] = 4'b1001;
	mem[3742] = 4'b1010;
	mem[3743] = 4'b1010;
	mem[3744] = 4'b1001;
	mem[3745] = 4'b1001;
	mem[3746] = 4'b1001;
	mem[3747] = 4'b0111;
	mem[3748] = 4'b0111;
	mem[3749] = 4'b0111;
	mem[3750] = 4'b0111;
	mem[3751] = 4'b0111;
	mem[3752] = 4'b1000;
	mem[3753] = 4'b0111;
	mem[3754] = 4'b0111;
	mem[3755] = 4'b0111;
	mem[3756] = 4'b0111;
	mem[3757] = 4'b0110;
	mem[3758] = 4'b0110;
	mem[3759] = 4'b0111;
	mem[3760] = 4'b0110;
	mem[3761] = 4'b0101;
	mem[3762] = 4'b0101;
	mem[3763] = 4'b0101;
	mem[3764] = 4'b0101;
	mem[3765] = 4'b0100;
	mem[3766] = 4'b0100;
	mem[3767] = 4'b0100;
	mem[3768] = 4'b0100;
	mem[3769] = 4'b0100;
	mem[3770] = 4'b0011;
	mem[3771] = 4'b0011;
	mem[3772] = 4'b0011;
	mem[3773] = 4'b0011;
	mem[3774] = 4'b0010;
	mem[3775] = 4'b0010;
	mem[3776] = 4'b0010;
	mem[3777] = 4'b0010;
	mem[3778] = 4'b0010;
	mem[3779] = 4'b0001;
	mem[3780] = 4'b0001;
	mem[3781] = 4'b0001;
	mem[3782] = 4'b0001;
	mem[3783] = 4'b0000;
	mem[3784] = 4'b0000;
	mem[3785] = 4'b0000;
	mem[3786] = 4'b0000;
	mem[3787] = 4'b1001;
	mem[3788] = 4'b1111;
	mem[3789] = 4'b1111;
	mem[3790] = 4'b1110;
	mem[3791] = 4'b1110;
	mem[3792] = 4'b1110;
	mem[3793] = 4'b1011;
	mem[3794] = 4'b1011;
	mem[3795] = 4'b1011;
	mem[3796] = 4'b1011;
	mem[3797] = 4'b1011;
	mem[3798] = 4'b1100;
	mem[3799] = 4'b1100;
	mem[3800] = 4'b1010;
	mem[3801] = 4'b1010;
	mem[3802] = 4'b1011;
	mem[3803] = 4'b1010;
	mem[3804] = 4'b1010;
	mem[3805] = 4'b1010;
	mem[3806] = 4'b1001;
	mem[3807] = 4'b1001;
	mem[3808] = 4'b1001;
	mem[3809] = 4'b1001;
	mem[3810] = 4'b1000;
	mem[3811] = 4'b1000;
	mem[3812] = 4'b1000;
	mem[3813] = 4'b1000;
	mem[3814] = 4'b0111;
	mem[3815] = 4'b0111;
	mem[3816] = 4'b0111;
	mem[3817] = 4'b0111;
	mem[3818] = 4'b0110;
	mem[3819] = 4'b0110;
	mem[3820] = 4'b0110;
	mem[3821] = 4'b0110;
	mem[3822] = 4'b0110;
	mem[3823] = 4'b0101;
	mem[3824] = 4'b0101;
	mem[3825] = 4'b0101;
	mem[3826] = 4'b0101;
	mem[3827] = 4'b0101;
	mem[3828] = 4'b0100;
	mem[3829] = 4'b0100;
	mem[3830] = 4'b0100;
	mem[3831] = 4'b0100;
	mem[3832] = 4'b0100;
	mem[3833] = 4'b0011;
	mem[3834] = 4'b0000;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b1001;
	mem[3844] = 4'b1111;
	mem[3845] = 4'b1111;
	mem[3846] = 4'b1111;
	mem[3847] = 4'b1111;
	mem[3848] = 4'b1110;
	mem[3849] = 4'b1110;
	mem[3850] = 4'b1110;
	mem[3851] = 4'b1110;
	mem[3852] = 4'b1101;
	mem[3853] = 4'b1101;
	mem[3854] = 4'b1101;
	mem[3855] = 4'b1101;
	mem[3856] = 4'b1101;
	mem[3857] = 4'b1100;
	mem[3858] = 4'b1100;
	mem[3859] = 4'b1100;
	mem[3860] = 4'b1100;
	mem[3861] = 4'b1011;
	mem[3862] = 4'b1011;
	mem[3863] = 4'b1011;
	mem[3864] = 4'b1011;
	mem[3865] = 4'b1010;
	mem[3866] = 4'b1001;
	mem[3867] = 4'b1001;
	mem[3868] = 4'b1001;
	mem[3869] = 4'b1010;
	mem[3870] = 4'b1010;
	mem[3871] = 4'b1001;
	mem[3872] = 4'b1001;
	mem[3873] = 4'b1001;
	mem[3874] = 4'b1001;
	mem[3875] = 4'b1001;
	mem[3876] = 4'b0111;
	mem[3877] = 4'b0111;
	mem[3878] = 4'b0111;
	mem[3879] = 4'b0111;
	mem[3880] = 4'b0111;
	mem[3881] = 4'b0111;
	mem[3882] = 4'b0111;
	mem[3883] = 4'b0111;
	mem[3884] = 4'b0110;
	mem[3885] = 4'b0111;
	mem[3886] = 4'b0111;
	mem[3887] = 4'b0110;
	mem[3888] = 4'b0101;
	mem[3889] = 4'b0101;
	mem[3890] = 4'b0101;
	mem[3891] = 4'b0101;
	mem[3892] = 4'b0101;
	mem[3893] = 4'b0100;
	mem[3894] = 4'b0100;
	mem[3895] = 4'b0100;
	mem[3896] = 4'b0100;
	mem[3897] = 4'b0100;
	mem[3898] = 4'b0011;
	mem[3899] = 4'b0011;
	mem[3900] = 4'b0011;
	mem[3901] = 4'b0011;
	mem[3902] = 4'b0010;
	mem[3903] = 4'b0010;
	mem[3904] = 4'b0010;
	mem[3905] = 4'b0010;
	mem[3906] = 4'b0010;
	mem[3907] = 4'b0001;
	mem[3908] = 4'b0001;
	mem[3909] = 4'b0001;
	mem[3910] = 4'b0001;
	mem[3911] = 4'b0000;
	mem[3912] = 4'b0000;
	mem[3913] = 4'b0000;
	mem[3914] = 4'b0000;
	mem[3915] = 4'b1001;
	mem[3916] = 4'b1111;
	mem[3917] = 4'b1110;
	mem[3918] = 4'b1110;
	mem[3919] = 4'b1110;
	mem[3920] = 4'b1110;
	mem[3921] = 4'b1101;
	mem[3922] = 4'b1100;
	mem[3923] = 4'b1100;
	mem[3924] = 4'b1100;
	mem[3925] = 4'b1100;
	mem[3926] = 4'b1100;
	mem[3927] = 4'b1011;
	mem[3928] = 4'b1010;
	mem[3929] = 4'b1011;
	mem[3930] = 4'b1011;
	mem[3931] = 4'b1010;
	mem[3932] = 4'b1010;
	mem[3933] = 4'b1010;
	mem[3934] = 4'b1001;
	mem[3935] = 4'b1001;
	mem[3936] = 4'b1001;
	mem[3937] = 4'b1001;
	mem[3938] = 4'b1000;
	mem[3939] = 4'b1000;
	mem[3940] = 4'b1000;
	mem[3941] = 4'b1000;
	mem[3942] = 4'b0111;
	mem[3943] = 4'b0111;
	mem[3944] = 4'b0111;
	mem[3945] = 4'b0111;
	mem[3946] = 4'b0111;
	mem[3947] = 4'b0110;
	mem[3948] = 4'b0110;
	mem[3949] = 4'b0110;
	mem[3950] = 4'b0110;
	mem[3951] = 4'b0110;
	mem[3952] = 4'b0101;
	mem[3953] = 4'b0101;
	mem[3954] = 4'b0101;
	mem[3955] = 4'b0101;
	mem[3956] = 4'b0101;
	mem[3957] = 4'b0100;
	mem[3958] = 4'b0100;
	mem[3959] = 4'b0100;
	mem[3960] = 4'b0100;
	mem[3961] = 4'b0100;
	mem[3962] = 4'b0001;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b1001;
	mem[3972] = 4'b1111;
	mem[3973] = 4'b1111;
	mem[3974] = 4'b1111;
	mem[3975] = 4'b1111;
	mem[3976] = 4'b1110;
	mem[3977] = 4'b1110;
	mem[3978] = 4'b1110;
	mem[3979] = 4'b1110;
	mem[3980] = 4'b1101;
	mem[3981] = 4'b1101;
	mem[3982] = 4'b1101;
	mem[3983] = 4'b1101;
	mem[3984] = 4'b1101;
	mem[3985] = 4'b1100;
	mem[3986] = 4'b1100;
	mem[3987] = 4'b1100;
	mem[3988] = 4'b1100;
	mem[3989] = 4'b1011;
	mem[3990] = 4'b1011;
	mem[3991] = 4'b1011;
	mem[3992] = 4'b1011;
	mem[3993] = 4'b1010;
	mem[3994] = 4'b1001;
	mem[3995] = 4'b1001;
	mem[3996] = 4'b1001;
	mem[3997] = 4'b1010;
	mem[3998] = 4'b1001;
	mem[3999] = 4'b1001;
	mem[4000] = 4'b1001;
	mem[4001] = 4'b1001;
	mem[4002] = 4'b1001;
	mem[4003] = 4'b1000;
	mem[4004] = 4'b1000;
	mem[4005] = 4'b0111;
	mem[4006] = 4'b0111;
	mem[4007] = 4'b0111;
	mem[4008] = 4'b0111;
	mem[4009] = 4'b0111;
	mem[4010] = 4'b0111;
	mem[4011] = 4'b0111;
	mem[4012] = 4'b0110;
	mem[4013] = 4'b0110;
	mem[4014] = 4'b0110;
	mem[4015] = 4'b0110;
	mem[4016] = 4'b0101;
	mem[4017] = 4'b0101;
	mem[4018] = 4'b0101;
	mem[4019] = 4'b0101;
	mem[4020] = 4'b0101;
	mem[4021] = 4'b0100;
	mem[4022] = 4'b0100;
	mem[4023] = 4'b0100;
	mem[4024] = 4'b0100;
	mem[4025] = 4'b0100;
	mem[4026] = 4'b0011;
	mem[4027] = 4'b0011;
	mem[4028] = 4'b0011;
	mem[4029] = 4'b0011;
	mem[4030] = 4'b0010;
	mem[4031] = 4'b0010;
	mem[4032] = 4'b0010;
	mem[4033] = 4'b0010;
	mem[4034] = 4'b0010;
	mem[4035] = 4'b0001;
	mem[4036] = 4'b0001;
	mem[4037] = 4'b0001;
	mem[4038] = 4'b0001;
	mem[4039] = 4'b0000;
	mem[4040] = 4'b0000;
	mem[4041] = 4'b0000;
	mem[4042] = 4'b0000;
	mem[4043] = 4'b1001;
	mem[4044] = 4'b1110;
	mem[4045] = 4'b1101;
	mem[4046] = 4'b1101;
	mem[4047] = 4'b1101;
	mem[4048] = 4'b1110;
	mem[4049] = 4'b1101;
	mem[4050] = 4'b1101;
	mem[4051] = 4'b1101;
	mem[4052] = 4'b1100;
	mem[4053] = 4'b1011;
	mem[4054] = 4'b1011;
	mem[4055] = 4'b1010;
	mem[4056] = 4'b1010;
	mem[4057] = 4'b1011;
	mem[4058] = 4'b1011;
	mem[4059] = 4'b1010;
	mem[4060] = 4'b1010;
	mem[4061] = 4'b1010;
	mem[4062] = 4'b1010;
	mem[4063] = 4'b1001;
	mem[4064] = 4'b1001;
	mem[4065] = 4'b1001;
	mem[4066] = 4'b1001;
	mem[4067] = 4'b1000;
	mem[4068] = 4'b1000;
	mem[4069] = 4'b1000;
	mem[4070] = 4'b1000;
	mem[4071] = 4'b0111;
	mem[4072] = 4'b0111;
	mem[4073] = 4'b0111;
	mem[4074] = 4'b0111;
	mem[4075] = 4'b0111;
	mem[4076] = 4'b0110;
	mem[4077] = 4'b0110;
	mem[4078] = 4'b0110;
	mem[4079] = 4'b0110;
	mem[4080] = 4'b0110;
	mem[4081] = 4'b0101;
	mem[4082] = 4'b0101;
	mem[4083] = 4'b0101;
	mem[4084] = 4'b0101;
	mem[4085] = 4'b0101;
	mem[4086] = 4'b0101;
	mem[4087] = 4'b0100;
	mem[4088] = 4'b0100;
	mem[4089] = 4'b0100;
	mem[4090] = 4'b0001;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_3r (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0110;
	mem[4] = 4'b1001;
	mem[5] = 4'b1001;
	mem[6] = 4'b1001;
	mem[7] = 4'b1001;
	mem[8] = 4'b1001;
	mem[9] = 4'b1001;
	mem[10] = 4'b1001;
	mem[11] = 4'b1001;
	mem[12] = 4'b1001;
	mem[13] = 4'b1001;
	mem[14] = 4'b1001;
	mem[15] = 4'b1001;
	mem[16] = 4'b1001;
	mem[17] = 4'b1001;
	mem[18] = 4'b1001;
	mem[19] = 4'b1000;
	mem[20] = 4'b1001;
	mem[21] = 4'b1001;
	mem[22] = 4'b1001;
	mem[23] = 4'b1001;
	mem[24] = 4'b1000;
	mem[25] = 4'b1000;
	mem[26] = 4'b1000;
	mem[27] = 4'b1000;
	mem[28] = 4'b1000;
	mem[29] = 4'b1001;
	mem[30] = 4'b1000;
	mem[31] = 4'b1000;
	mem[32] = 4'b1000;
	mem[33] = 4'b1000;
	mem[34] = 4'b1000;
	mem[35] = 4'b1000;
	mem[36] = 4'b1000;
	mem[37] = 4'b1000;
	mem[38] = 4'b0111;
	mem[39] = 4'b0111;
	mem[40] = 4'b0111;
	mem[41] = 4'b1000;
	mem[42] = 4'b1000;
	mem[43] = 4'b1000;
	mem[44] = 4'b1000;
	mem[45] = 4'b1000;
	mem[46] = 4'b1000;
	mem[47] = 4'b1000;
	mem[48] = 4'b1000;
	mem[49] = 4'b1000;
	mem[50] = 4'b1000;
	mem[51] = 4'b1000;
	mem[52] = 4'b0111;
	mem[53] = 4'b1000;
	mem[54] = 4'b1000;
	mem[55] = 4'b1000;
	mem[56] = 4'b1000;
	mem[57] = 4'b0111;
	mem[58] = 4'b0111;
	mem[59] = 4'b0111;
	mem[60] = 4'b0111;
	mem[61] = 4'b0111;
	mem[62] = 4'b0111;
	mem[63] = 4'b0111;
	mem[64] = 4'b0111;
	mem[65] = 4'b0111;
	mem[66] = 4'b0111;
	mem[67] = 4'b0111;
	mem[68] = 4'b0111;
	mem[69] = 4'b0110;
	mem[70] = 4'b0011;
	mem[71] = 4'b0000;
	mem[72] = 4'b0000;
	mem[73] = 4'b0000;
	mem[74] = 4'b0000;
	mem[75] = 4'b0101;
	mem[76] = 4'b1000;
	mem[77] = 4'b1000;
	mem[78] = 4'b1000;
	mem[79] = 4'b1000;
	mem[80] = 4'b1000;
	mem[81] = 4'b1000;
	mem[82] = 4'b1000;
	mem[83] = 4'b1000;
	mem[84] = 4'b0111;
	mem[85] = 4'b0111;
	mem[86] = 4'b0111;
	mem[87] = 4'b1000;
	mem[88] = 4'b1000;
	mem[89] = 4'b0111;
	mem[90] = 4'b0111;
	mem[91] = 4'b0111;
	mem[92] = 4'b0111;
	mem[93] = 4'b0111;
	mem[94] = 4'b0111;
	mem[95] = 4'b0110;
	mem[96] = 4'b0110;
	mem[97] = 4'b0110;
	mem[98] = 4'b0110;
	mem[99] = 4'b0110;
	mem[100] = 4'b0110;
	mem[101] = 4'b0110;
	mem[102] = 4'b0110;
	mem[103] = 4'b0110;
	mem[104] = 4'b0101;
	mem[105] = 4'b0101;
	mem[106] = 4'b0101;
	mem[107] = 4'b0101;
	mem[108] = 4'b0101;
	mem[109] = 4'b0101;
	mem[110] = 4'b0101;
	mem[111] = 4'b0101;
	mem[112] = 4'b0101;
	mem[113] = 4'b0101;
	mem[114] = 4'b0101;
	mem[115] = 4'b0101;
	mem[116] = 4'b0101;
	mem[117] = 4'b0101;
	mem[118] = 4'b0101;
	mem[119] = 4'b0100;
	mem[120] = 4'b0100;
	mem[121] = 4'b0100;
	mem[122] = 4'b0001;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b0000;
	mem[132] = 4'b0000;
	mem[133] = 4'b0000;
	mem[134] = 4'b0000;
	mem[135] = 4'b0000;
	mem[136] = 4'b0000;
	mem[137] = 4'b0001;
	mem[138] = 4'b0001;
	mem[139] = 4'b0001;
	mem[140] = 4'b0001;
	mem[141] = 4'b0001;
	mem[142] = 4'b0010;
	mem[143] = 4'b0011;
	mem[144] = 4'b0011;
	mem[145] = 4'b0011;
	mem[146] = 4'b0011;
	mem[147] = 4'b0011;
	mem[148] = 4'b0100;
	mem[149] = 4'b0100;
	mem[150] = 4'b0100;
	mem[151] = 4'b0100;
	mem[152] = 4'b0100;
	mem[153] = 4'b0101;
	mem[154] = 4'b0101;
	mem[155] = 4'b0101;
	mem[156] = 4'b0110;
	mem[157] = 4'b0110;
	mem[158] = 4'b0110;
	mem[159] = 4'b0111;
	mem[160] = 4'b1000;
	mem[161] = 4'b1000;
	mem[162] = 4'b1000;
	mem[163] = 4'b1000;
	mem[164] = 4'b1000;
	mem[165] = 4'b1001;
	mem[166] = 4'b1000;
	mem[167] = 4'b1000;
	mem[168] = 4'b1000;
	mem[169] = 4'b1001;
	mem[170] = 4'b1010;
	mem[171] = 4'b1011;
	mem[172] = 4'b1011;
	mem[173] = 4'b1011;
	mem[174] = 4'b1011;
	mem[175] = 4'b1011;
	mem[176] = 4'b1100;
	mem[177] = 4'b1100;
	mem[178] = 4'b1100;
	mem[179] = 4'b1100;
	mem[180] = 4'b1100;
	mem[181] = 4'b1101;
	mem[182] = 4'b1110;
	mem[183] = 4'b1110;
	mem[184] = 4'b1110;
	mem[185] = 4'b1110;
	mem[186] = 4'b1110;
	mem[187] = 4'b1111;
	mem[188] = 4'b1111;
	mem[189] = 4'b1111;
	mem[190] = 4'b1111;
	mem[191] = 4'b1111;
	mem[192] = 4'b1111;
	mem[193] = 4'b1111;
	mem[194] = 4'b1111;
	mem[195] = 4'b1111;
	mem[196] = 4'b1111;
	mem[197] = 4'b1111;
	mem[198] = 4'b0110;
	mem[199] = 4'b0000;
	mem[200] = 4'b0000;
	mem[201] = 4'b0000;
	mem[202] = 4'b0000;
	mem[203] = 4'b0000;
	mem[204] = 4'b0001;
	mem[205] = 4'b0001;
	mem[206] = 4'b0001;
	mem[207] = 4'b0000;
	mem[208] = 4'b0000;
	mem[209] = 4'b0001;
	mem[210] = 4'b0001;
	mem[211] = 4'b0000;
	mem[212] = 4'b0001;
	mem[213] = 4'b0010;
	mem[214] = 4'b0010;
	mem[215] = 4'b0010;
	mem[216] = 4'b0001;
	mem[217] = 4'b0001;
	mem[218] = 4'b0001;
	mem[219] = 4'b0001;
	mem[220] = 4'b0001;
	mem[221] = 4'b0001;
	mem[222] = 4'b0010;
	mem[223] = 4'b0010;
	mem[224] = 4'b0010;
	mem[225] = 4'b0010;
	mem[226] = 4'b0010;
	mem[227] = 4'b0010;
	mem[228] = 4'b0010;
	mem[229] = 4'b0010;
	mem[230] = 4'b0010;
	mem[231] = 4'b0011;
	mem[232] = 4'b0011;
	mem[233] = 4'b0011;
	mem[234] = 4'b0011;
	mem[235] = 4'b0011;
	mem[236] = 4'b0011;
	mem[237] = 4'b0011;
	mem[238] = 4'b0011;
	mem[239] = 4'b0011;
	mem[240] = 4'b0100;
	mem[241] = 4'b0100;
	mem[242] = 4'b0100;
	mem[243] = 4'b0100;
	mem[244] = 4'b0100;
	mem[245] = 4'b0100;
	mem[246] = 4'b0100;
	mem[247] = 4'b0100;
	mem[248] = 4'b0100;
	mem[249] = 4'b0100;
	mem[250] = 4'b0001;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0000;
	mem[260] = 4'b0000;
	mem[261] = 4'b0000;
	mem[262] = 4'b0000;
	mem[263] = 4'b0000;
	mem[264] = 4'b0000;
	mem[265] = 4'b0001;
	mem[266] = 4'b0001;
	mem[267] = 4'b0001;
	mem[268] = 4'b0001;
	mem[269] = 4'b0001;
	mem[270] = 4'b0010;
	mem[271] = 4'b0011;
	mem[272] = 4'b0011;
	mem[273] = 4'b0011;
	mem[274] = 4'b0011;
	mem[275] = 4'b0011;
	mem[276] = 4'b0100;
	mem[277] = 4'b0100;
	mem[278] = 4'b0100;
	mem[279] = 4'b0100;
	mem[280] = 4'b0100;
	mem[281] = 4'b0101;
	mem[282] = 4'b0101;
	mem[283] = 4'b0101;
	mem[284] = 4'b0101;
	mem[285] = 4'b0110;
	mem[286] = 4'b0110;
	mem[287] = 4'b0111;
	mem[288] = 4'b1000;
	mem[289] = 4'b1000;
	mem[290] = 4'b1000;
	mem[291] = 4'b1000;
	mem[292] = 4'b1000;
	mem[293] = 4'b1000;
	mem[294] = 4'b1000;
	mem[295] = 4'b1000;
	mem[296] = 4'b1001;
	mem[297] = 4'b1001;
	mem[298] = 4'b1010;
	mem[299] = 4'b1011;
	mem[300] = 4'b1011;
	mem[301] = 4'b1011;
	mem[302] = 4'b1011;
	mem[303] = 4'b1011;
	mem[304] = 4'b1100;
	mem[305] = 4'b1100;
	mem[306] = 4'b1100;
	mem[307] = 4'b1100;
	mem[308] = 4'b1100;
	mem[309] = 4'b1101;
	mem[310] = 4'b1110;
	mem[311] = 4'b1110;
	mem[312] = 4'b1110;
	mem[313] = 4'b1110;
	mem[314] = 4'b1110;
	mem[315] = 4'b1111;
	mem[316] = 4'b1111;
	mem[317] = 4'b1111;
	mem[318] = 4'b1111;
	mem[319] = 4'b1111;
	mem[320] = 4'b1111;
	mem[321] = 4'b1111;
	mem[322] = 4'b1111;
	mem[323] = 4'b1111;
	mem[324] = 4'b1111;
	mem[325] = 4'b1111;
	mem[326] = 4'b0110;
	mem[327] = 4'b0000;
	mem[328] = 4'b0000;
	mem[329] = 4'b0000;
	mem[330] = 4'b0000;
	mem[331] = 4'b0000;
	mem[332] = 4'b0001;
	mem[333] = 4'b0000;
	mem[334] = 4'b0000;
	mem[335] = 4'b0001;
	mem[336] = 4'b0001;
	mem[337] = 4'b0001;
	mem[338] = 4'b0001;
	mem[339] = 4'b0001;
	mem[340] = 4'b0001;
	mem[341] = 4'b0001;
	mem[342] = 4'b0001;
	mem[343] = 4'b0001;
	mem[344] = 4'b0001;
	mem[345] = 4'b0001;
	mem[346] = 4'b0001;
	mem[347] = 4'b0010;
	mem[348] = 4'b0010;
	mem[349] = 4'b0010;
	mem[350] = 4'b0010;
	mem[351] = 4'b0010;
	mem[352] = 4'b0010;
	mem[353] = 4'b0010;
	mem[354] = 4'b0010;
	mem[355] = 4'b0010;
	mem[356] = 4'b0011;
	mem[357] = 4'b0011;
	mem[358] = 4'b0011;
	mem[359] = 4'b0011;
	mem[360] = 4'b0011;
	mem[361] = 4'b0011;
	mem[362] = 4'b0011;
	mem[363] = 4'b0011;
	mem[364] = 4'b0011;
	mem[365] = 4'b0011;
	mem[366] = 4'b0100;
	mem[367] = 4'b0100;
	mem[368] = 4'b0100;
	mem[369] = 4'b0100;
	mem[370] = 4'b0100;
	mem[371] = 4'b0100;
	mem[372] = 4'b0100;
	mem[373] = 4'b0100;
	mem[374] = 4'b0100;
	mem[375] = 4'b0101;
	mem[376] = 4'b0101;
	mem[377] = 4'b0101;
	mem[378] = 4'b0001;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0000;
	mem[388] = 4'b0000;
	mem[389] = 4'b0000;
	mem[390] = 4'b0000;
	mem[391] = 4'b0000;
	mem[392] = 4'b0000;
	mem[393] = 4'b0001;
	mem[394] = 4'b0001;
	mem[395] = 4'b0001;
	mem[396] = 4'b0001;
	mem[397] = 4'b0001;
	mem[398] = 4'b0010;
	mem[399] = 4'b0011;
	mem[400] = 4'b0011;
	mem[401] = 4'b0011;
	mem[402] = 4'b0011;
	mem[403] = 4'b0011;
	mem[404] = 4'b0100;
	mem[405] = 4'b0100;
	mem[406] = 4'b0100;
	mem[407] = 4'b0100;
	mem[408] = 4'b0100;
	mem[409] = 4'b0101;
	mem[410] = 4'b0101;
	mem[411] = 4'b0101;
	mem[412] = 4'b0101;
	mem[413] = 4'b0101;
	mem[414] = 4'b0110;
	mem[415] = 4'b0111;
	mem[416] = 4'b1000;
	mem[417] = 4'b1000;
	mem[418] = 4'b1000;
	mem[419] = 4'b1000;
	mem[420] = 4'b1000;
	mem[421] = 4'b1000;
	mem[422] = 4'b1000;
	mem[423] = 4'b1000;
	mem[424] = 4'b1001;
	mem[425] = 4'b1001;
	mem[426] = 4'b1010;
	mem[427] = 4'b1011;
	mem[428] = 4'b1011;
	mem[429] = 4'b1011;
	mem[430] = 4'b1011;
	mem[431] = 4'b1011;
	mem[432] = 4'b1100;
	mem[433] = 4'b1100;
	mem[434] = 4'b1100;
	mem[435] = 4'b1100;
	mem[436] = 4'b1100;
	mem[437] = 4'b1101;
	mem[438] = 4'b1110;
	mem[439] = 4'b1110;
	mem[440] = 4'b1110;
	mem[441] = 4'b1110;
	mem[442] = 4'b1110;
	mem[443] = 4'b1111;
	mem[444] = 4'b1111;
	mem[445] = 4'b1111;
	mem[446] = 4'b1111;
	mem[447] = 4'b1111;
	mem[448] = 4'b1111;
	mem[449] = 4'b1111;
	mem[450] = 4'b1111;
	mem[451] = 4'b1111;
	mem[452] = 4'b1111;
	mem[453] = 4'b1111;
	mem[454] = 4'b0110;
	mem[455] = 4'b0000;
	mem[456] = 4'b0000;
	mem[457] = 4'b0000;
	mem[458] = 4'b0000;
	mem[459] = 4'b0001;
	mem[460] = 4'b0001;
	mem[461] = 4'b0000;
	mem[462] = 4'b0000;
	mem[463] = 4'b0001;
	mem[464] = 4'b0001;
	mem[465] = 4'b0001;
	mem[466] = 4'b0001;
	mem[467] = 4'b0010;
	mem[468] = 4'b0001;
	mem[469] = 4'b0001;
	mem[470] = 4'b0001;
	mem[471] = 4'b0001;
	mem[472] = 4'b0001;
	mem[473] = 4'b0010;
	mem[474] = 4'b0010;
	mem[475] = 4'b0010;
	mem[476] = 4'b0010;
	mem[477] = 4'b0010;
	mem[478] = 4'b0010;
	mem[479] = 4'b0010;
	mem[480] = 4'b0010;
	mem[481] = 4'b0010;
	mem[482] = 4'b0011;
	mem[483] = 4'b0011;
	mem[484] = 4'b0011;
	mem[485] = 4'b0011;
	mem[486] = 4'b0011;
	mem[487] = 4'b0011;
	mem[488] = 4'b0011;
	mem[489] = 4'b0011;
	mem[490] = 4'b0011;
	mem[491] = 4'b0100;
	mem[492] = 4'b0100;
	mem[493] = 4'b0100;
	mem[494] = 4'b0100;
	mem[495] = 4'b0100;
	mem[496] = 4'b0100;
	mem[497] = 4'b0100;
	mem[498] = 4'b0100;
	mem[499] = 4'b0100;
	mem[500] = 4'b0101;
	mem[501] = 4'b0101;
	mem[502] = 4'b0101;
	mem[503] = 4'b0101;
	mem[504] = 4'b0101;
	mem[505] = 4'b0101;
	mem[506] = 4'b0001;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0000;
	mem[516] = 4'b0000;
	mem[517] = 4'b0000;
	mem[518] = 4'b0000;
	mem[519] = 4'b0000;
	mem[520] = 4'b0000;
	mem[521] = 4'b0001;
	mem[522] = 4'b0001;
	mem[523] = 4'b0001;
	mem[524] = 4'b0001;
	mem[525] = 4'b0001;
	mem[526] = 4'b0010;
	mem[527] = 4'b0011;
	mem[528] = 4'b0011;
	mem[529] = 4'b0011;
	mem[530] = 4'b0011;
	mem[531] = 4'b0011;
	mem[532] = 4'b0100;
	mem[533] = 4'b0100;
	mem[534] = 4'b0100;
	mem[535] = 4'b0100;
	mem[536] = 4'b0100;
	mem[537] = 4'b0101;
	mem[538] = 4'b0110;
	mem[539] = 4'b0101;
	mem[540] = 4'b0101;
	mem[541] = 4'b0101;
	mem[542] = 4'b0101;
	mem[543] = 4'b0111;
	mem[544] = 4'b1000;
	mem[545] = 4'b1000;
	mem[546] = 4'b0111;
	mem[547] = 4'b0111;
	mem[548] = 4'b0111;
	mem[549] = 4'b1000;
	mem[550] = 4'b1000;
	mem[551] = 4'b1000;
	mem[552] = 4'b1010;
	mem[553] = 4'b1001;
	mem[554] = 4'b1010;
	mem[555] = 4'b1011;
	mem[556] = 4'b1011;
	mem[557] = 4'b1011;
	mem[558] = 4'b1011;
	mem[559] = 4'b1011;
	mem[560] = 4'b1100;
	mem[561] = 4'b1100;
	mem[562] = 4'b1100;
	mem[563] = 4'b1100;
	mem[564] = 4'b1100;
	mem[565] = 4'b1101;
	mem[566] = 4'b1110;
	mem[567] = 4'b1110;
	mem[568] = 4'b1110;
	mem[569] = 4'b1110;
	mem[570] = 4'b1110;
	mem[571] = 4'b1111;
	mem[572] = 4'b1111;
	mem[573] = 4'b1111;
	mem[574] = 4'b1111;
	mem[575] = 4'b1111;
	mem[576] = 4'b1111;
	mem[577] = 4'b1111;
	mem[578] = 4'b1111;
	mem[579] = 4'b1111;
	mem[580] = 4'b1111;
	mem[581] = 4'b1111;
	mem[582] = 4'b0110;
	mem[583] = 4'b0000;
	mem[584] = 4'b0000;
	mem[585] = 4'b0001;
	mem[586] = 4'b0001;
	mem[587] = 4'b0001;
	mem[588] = 4'b0001;
	mem[589] = 4'b0001;
	mem[590] = 4'b0001;
	mem[591] = 4'b0001;
	mem[592] = 4'b0001;
	mem[593] = 4'b0010;
	mem[594] = 4'b0001;
	mem[595] = 4'b0010;
	mem[596] = 4'b0010;
	mem[597] = 4'b0001;
	mem[598] = 4'b0010;
	mem[599] = 4'b0010;
	mem[600] = 4'b0010;
	mem[601] = 4'b0010;
	mem[602] = 4'b0010;
	mem[603] = 4'b0010;
	mem[604] = 4'b0010;
	mem[605] = 4'b0010;
	mem[606] = 4'b0010;
	mem[607] = 4'b0011;
	mem[608] = 4'b0011;
	mem[609] = 4'b0011;
	mem[610] = 4'b0011;
	mem[611] = 4'b0011;
	mem[612] = 4'b0011;
	mem[613] = 4'b0011;
	mem[614] = 4'b0011;
	mem[615] = 4'b0011;
	mem[616] = 4'b0100;
	mem[617] = 4'b0100;
	mem[618] = 4'b0100;
	mem[619] = 4'b0100;
	mem[620] = 4'b0100;
	mem[621] = 4'b0100;
	mem[622] = 4'b0100;
	mem[623] = 4'b0100;
	mem[624] = 4'b0100;
	mem[625] = 4'b0100;
	mem[626] = 4'b0101;
	mem[627] = 4'b0101;
	mem[628] = 4'b0101;
	mem[629] = 4'b0101;
	mem[630] = 4'b0101;
	mem[631] = 4'b0101;
	mem[632] = 4'b0101;
	mem[633] = 4'b0101;
	mem[634] = 4'b0001;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0000;
	mem[644] = 4'b0000;
	mem[645] = 4'b0000;
	mem[646] = 4'b0000;
	mem[647] = 4'b0000;
	mem[648] = 4'b0000;
	mem[649] = 4'b0001;
	mem[650] = 4'b0001;
	mem[651] = 4'b0001;
	mem[652] = 4'b0001;
	mem[653] = 4'b0001;
	mem[654] = 4'b0010;
	mem[655] = 4'b0011;
	mem[656] = 4'b0011;
	mem[657] = 4'b0011;
	mem[658] = 4'b0011;
	mem[659] = 4'b0011;
	mem[660] = 4'b0100;
	mem[661] = 4'b0100;
	mem[662] = 4'b0100;
	mem[663] = 4'b0101;
	mem[664] = 4'b0100;
	mem[665] = 4'b0101;
	mem[666] = 4'b0110;
	mem[667] = 4'b0101;
	mem[668] = 4'b0101;
	mem[669] = 4'b0101;
	mem[670] = 4'b0101;
	mem[671] = 4'b0110;
	mem[672] = 4'b0111;
	mem[673] = 4'b0111;
	mem[674] = 4'b0111;
	mem[675] = 4'b0111;
	mem[676] = 4'b0111;
	mem[677] = 4'b1000;
	mem[678] = 4'b1000;
	mem[679] = 4'b1001;
	mem[680] = 4'b1001;
	mem[681] = 4'b1001;
	mem[682] = 4'b1010;
	mem[683] = 4'b1011;
	mem[684] = 4'b1011;
	mem[685] = 4'b1011;
	mem[686] = 4'b1011;
	mem[687] = 4'b1011;
	mem[688] = 4'b1100;
	mem[689] = 4'b1100;
	mem[690] = 4'b1100;
	mem[691] = 4'b1100;
	mem[692] = 4'b1100;
	mem[693] = 4'b1101;
	mem[694] = 4'b1110;
	mem[695] = 4'b1110;
	mem[696] = 4'b1110;
	mem[697] = 4'b1110;
	mem[698] = 4'b1110;
	mem[699] = 4'b1111;
	mem[700] = 4'b1111;
	mem[701] = 4'b1111;
	mem[702] = 4'b1111;
	mem[703] = 4'b1111;
	mem[704] = 4'b1111;
	mem[705] = 4'b1111;
	mem[706] = 4'b1111;
	mem[707] = 4'b1111;
	mem[708] = 4'b1111;
	mem[709] = 4'b1111;
	mem[710] = 4'b0110;
	mem[711] = 4'b0000;
	mem[712] = 4'b0000;
	mem[713] = 4'b0000;
	mem[714] = 4'b0001;
	mem[715] = 4'b0001;
	mem[716] = 4'b0001;
	mem[717] = 4'b0010;
	mem[718] = 4'b0001;
	mem[719] = 4'b0001;
	mem[720] = 4'b0001;
	mem[721] = 4'b0001;
	mem[722] = 4'b0010;
	mem[723] = 4'b0011;
	mem[724] = 4'b0010;
	mem[725] = 4'b0010;
	mem[726] = 4'b0010;
	mem[727] = 4'b0010;
	mem[728] = 4'b0010;
	mem[729] = 4'b0010;
	mem[730] = 4'b0010;
	mem[731] = 4'b0010;
	mem[732] = 4'b0010;
	mem[733] = 4'b0011;
	mem[734] = 4'b0011;
	mem[735] = 4'b0011;
	mem[736] = 4'b0011;
	mem[737] = 4'b0011;
	mem[738] = 4'b0011;
	mem[739] = 4'b0011;
	mem[740] = 4'b0011;
	mem[741] = 4'b0011;
	mem[742] = 4'b0100;
	mem[743] = 4'b0100;
	mem[744] = 4'b0100;
	mem[745] = 4'b0100;
	mem[746] = 4'b0100;
	mem[747] = 4'b0100;
	mem[748] = 4'b0100;
	mem[749] = 4'b0100;
	mem[750] = 4'b0100;
	mem[751] = 4'b0101;
	mem[752] = 4'b0101;
	mem[753] = 4'b0101;
	mem[754] = 4'b0101;
	mem[755] = 4'b0101;
	mem[756] = 4'b0101;
	mem[757] = 4'b0101;
	mem[758] = 4'b0101;
	mem[759] = 4'b0101;
	mem[760] = 4'b0110;
	mem[761] = 4'b0101;
	mem[762] = 4'b0001;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0000;
	mem[772] = 4'b0000;
	mem[773] = 4'b0000;
	mem[774] = 4'b0000;
	mem[775] = 4'b0000;
	mem[776] = 4'b0000;
	mem[777] = 4'b0001;
	mem[778] = 4'b0001;
	mem[779] = 4'b0001;
	mem[780] = 4'b0001;
	mem[781] = 4'b0001;
	mem[782] = 4'b0010;
	mem[783] = 4'b0011;
	mem[784] = 4'b0011;
	mem[785] = 4'b0011;
	mem[786] = 4'b0011;
	mem[787] = 4'b0011;
	mem[788] = 4'b0100;
	mem[789] = 4'b0100;
	mem[790] = 4'b0100;
	mem[791] = 4'b0101;
	mem[792] = 4'b0101;
	mem[793] = 4'b0101;
	mem[794] = 4'b0110;
	mem[795] = 4'b0110;
	mem[796] = 4'b0101;
	mem[797] = 4'b0101;
	mem[798] = 4'b0101;
	mem[799] = 4'b0110;
	mem[800] = 4'b0111;
	mem[801] = 4'b0111;
	mem[802] = 4'b0111;
	mem[803] = 4'b0111;
	mem[804] = 4'b0111;
	mem[805] = 4'b1000;
	mem[806] = 4'b1001;
	mem[807] = 4'b1010;
	mem[808] = 4'b1001;
	mem[809] = 4'b1001;
	mem[810] = 4'b1010;
	mem[811] = 4'b1011;
	mem[812] = 4'b1011;
	mem[813] = 4'b1011;
	mem[814] = 4'b1011;
	mem[815] = 4'b1011;
	mem[816] = 4'b1100;
	mem[817] = 4'b1100;
	mem[818] = 4'b1100;
	mem[819] = 4'b1100;
	mem[820] = 4'b1100;
	mem[821] = 4'b1101;
	mem[822] = 4'b1110;
	mem[823] = 4'b1110;
	mem[824] = 4'b1110;
	mem[825] = 4'b1110;
	mem[826] = 4'b1110;
	mem[827] = 4'b1111;
	mem[828] = 4'b1111;
	mem[829] = 4'b1111;
	mem[830] = 4'b1111;
	mem[831] = 4'b1111;
	mem[832] = 4'b1111;
	mem[833] = 4'b1111;
	mem[834] = 4'b1111;
	mem[835] = 4'b1111;
	mem[836] = 4'b1111;
	mem[837] = 4'b1110;
	mem[838] = 4'b0110;
	mem[839] = 4'b0001;
	mem[840] = 4'b0001;
	mem[841] = 4'b0001;
	mem[842] = 4'b0001;
	mem[843] = 4'b0010;
	mem[844] = 4'b0001;
	mem[845] = 4'b0001;
	mem[846] = 4'b0010;
	mem[847] = 4'b0010;
	mem[848] = 4'b0001;
	mem[849] = 4'b0010;
	mem[850] = 4'b0010;
	mem[851] = 4'b0010;
	mem[852] = 4'b0010;
	mem[853] = 4'b0010;
	mem[854] = 4'b0010;
	mem[855] = 4'b0010;
	mem[856] = 4'b0010;
	mem[857] = 4'b0010;
	mem[858] = 4'b0011;
	mem[859] = 4'b0011;
	mem[860] = 4'b0011;
	mem[861] = 4'b0011;
	mem[862] = 4'b0011;
	mem[863] = 4'b0011;
	mem[864] = 4'b0011;
	mem[865] = 4'b0011;
	mem[866] = 4'b0011;
	mem[867] = 4'b0100;
	mem[868] = 4'b0100;
	mem[869] = 4'b0100;
	mem[870] = 4'b0100;
	mem[871] = 4'b0100;
	mem[872] = 4'b0100;
	mem[873] = 4'b0100;
	mem[874] = 4'b0100;
	mem[875] = 4'b0100;
	mem[876] = 4'b0101;
	mem[877] = 4'b0101;
	mem[878] = 4'b0101;
	mem[879] = 4'b0101;
	mem[880] = 4'b0101;
	mem[881] = 4'b0101;
	mem[882] = 4'b0101;
	mem[883] = 4'b0101;
	mem[884] = 4'b0101;
	mem[885] = 4'b0101;
	mem[886] = 4'b0110;
	mem[887] = 4'b0110;
	mem[888] = 4'b0110;
	mem[889] = 4'b0110;
	mem[890] = 4'b0001;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0000;
	mem[900] = 4'b0000;
	mem[901] = 4'b0000;
	mem[902] = 4'b0000;
	mem[903] = 4'b0000;
	mem[904] = 4'b0000;
	mem[905] = 4'b0001;
	mem[906] = 4'b0001;
	mem[907] = 4'b0001;
	mem[908] = 4'b0001;
	mem[909] = 4'b0001;
	mem[910] = 4'b0010;
	mem[911] = 4'b0011;
	mem[912] = 4'b0011;
	mem[913] = 4'b0011;
	mem[914] = 4'b0011;
	mem[915] = 4'b0011;
	mem[916] = 4'b0100;
	mem[917] = 4'b0100;
	mem[918] = 4'b0101;
	mem[919] = 4'b0101;
	mem[920] = 4'b0100;
	mem[921] = 4'b0101;
	mem[922] = 4'b0110;
	mem[923] = 4'b0110;
	mem[924] = 4'b0110;
	mem[925] = 4'b0110;
	mem[926] = 4'b0101;
	mem[927] = 4'b0110;
	mem[928] = 4'b0111;
	mem[929] = 4'b0111;
	mem[930] = 4'b0111;
	mem[931] = 4'b0111;
	mem[932] = 4'b0111;
	mem[933] = 4'b1001;
	mem[934] = 4'b1010;
	mem[935] = 4'b1001;
	mem[936] = 4'b1001;
	mem[937] = 4'b1001;
	mem[938] = 4'b1010;
	mem[939] = 4'b1011;
	mem[940] = 4'b1011;
	mem[941] = 4'b1011;
	mem[942] = 4'b1011;
	mem[943] = 4'b1011;
	mem[944] = 4'b1100;
	mem[945] = 4'b1100;
	mem[946] = 4'b1100;
	mem[947] = 4'b1100;
	mem[948] = 4'b1100;
	mem[949] = 4'b1101;
	mem[950] = 4'b1110;
	mem[951] = 4'b1110;
	mem[952] = 4'b1110;
	mem[953] = 4'b1110;
	mem[954] = 4'b1110;
	mem[955] = 4'b1111;
	mem[956] = 4'b1111;
	mem[957] = 4'b1111;
	mem[958] = 4'b1111;
	mem[959] = 4'b1111;
	mem[960] = 4'b1111;
	mem[961] = 4'b1111;
	mem[962] = 4'b1111;
	mem[963] = 4'b1111;
	mem[964] = 4'b1110;
	mem[965] = 4'b1101;
	mem[966] = 4'b0110;
	mem[967] = 4'b0001;
	mem[968] = 4'b0001;
	mem[969] = 4'b0001;
	mem[970] = 4'b0010;
	mem[971] = 4'b0001;
	mem[972] = 4'b0010;
	mem[973] = 4'b0010;
	mem[974] = 4'b0010;
	mem[975] = 4'b0010;
	mem[976] = 4'b0010;
	mem[977] = 4'b0010;
	mem[978] = 4'b0010;
	mem[979] = 4'b0010;
	mem[980] = 4'b0010;
	mem[981] = 4'b0010;
	mem[982] = 4'b0010;
	mem[983] = 4'b0010;
	mem[984] = 4'b0011;
	mem[985] = 4'b0011;
	mem[986] = 4'b0011;
	mem[987] = 4'b0011;
	mem[988] = 4'b0011;
	mem[989] = 4'b0011;
	mem[990] = 4'b0011;
	mem[991] = 4'b0011;
	mem[992] = 4'b0011;
	mem[993] = 4'b0100;
	mem[994] = 4'b0100;
	mem[995] = 4'b0100;
	mem[996] = 4'b0100;
	mem[997] = 4'b0100;
	mem[998] = 4'b0100;
	mem[999] = 4'b0100;
	mem[1000] = 4'b0100;
	mem[1001] = 4'b0100;
	mem[1002] = 4'b0101;
	mem[1003] = 4'b0101;
	mem[1004] = 4'b0101;
	mem[1005] = 4'b0101;
	mem[1006] = 4'b0101;
	mem[1007] = 4'b0101;
	mem[1008] = 4'b0101;
	mem[1009] = 4'b0101;
	mem[1010] = 4'b0101;
	mem[1011] = 4'b0110;
	mem[1012] = 4'b0110;
	mem[1013] = 4'b0110;
	mem[1014] = 4'b0110;
	mem[1015] = 4'b0110;
	mem[1016] = 4'b0110;
	mem[1017] = 4'b0110;
	mem[1018] = 4'b0001;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0000;
	mem[1028] = 4'b0000;
	mem[1029] = 4'b0000;
	mem[1030] = 4'b0000;
	mem[1031] = 4'b0000;
	mem[1032] = 4'b0000;
	mem[1033] = 4'b0001;
	mem[1034] = 4'b0001;
	mem[1035] = 4'b0001;
	mem[1036] = 4'b0001;
	mem[1037] = 4'b0001;
	mem[1038] = 4'b0010;
	mem[1039] = 4'b0011;
	mem[1040] = 4'b0011;
	mem[1041] = 4'b0011;
	mem[1042] = 4'b0011;
	mem[1043] = 4'b0100;
	mem[1044] = 4'b0101;
	mem[1045] = 4'b0101;
	mem[1046] = 4'b0101;
	mem[1047] = 4'b0100;
	mem[1048] = 4'b0100;
	mem[1049] = 4'b0101;
	mem[1050] = 4'b0110;
	mem[1051] = 4'b0110;
	mem[1052] = 4'b0110;
	mem[1053] = 4'b0110;
	mem[1054] = 4'b0110;
	mem[1055] = 4'b0111;
	mem[1056] = 4'b0111;
	mem[1057] = 4'b0111;
	mem[1058] = 4'b0111;
	mem[1059] = 4'b1000;
	mem[1060] = 4'b1000;
	mem[1061] = 4'b1001;
	mem[1062] = 4'b1001;
	mem[1063] = 4'b1001;
	mem[1064] = 4'b1001;
	mem[1065] = 4'b1001;
	mem[1066] = 4'b1010;
	mem[1067] = 4'b1011;
	mem[1068] = 4'b1011;
	mem[1069] = 4'b1011;
	mem[1070] = 4'b1011;
	mem[1071] = 4'b1011;
	mem[1072] = 4'b1100;
	mem[1073] = 4'b1100;
	mem[1074] = 4'b1100;
	mem[1075] = 4'b1100;
	mem[1076] = 4'b1100;
	mem[1077] = 4'b1101;
	mem[1078] = 4'b1110;
	mem[1079] = 4'b1110;
	mem[1080] = 4'b1110;
	mem[1081] = 4'b1110;
	mem[1082] = 4'b1110;
	mem[1083] = 4'b1111;
	mem[1084] = 4'b1111;
	mem[1085] = 4'b1111;
	mem[1086] = 4'b1111;
	mem[1087] = 4'b1111;
	mem[1088] = 4'b1111;
	mem[1089] = 4'b1111;
	mem[1090] = 4'b1111;
	mem[1091] = 4'b1110;
	mem[1092] = 4'b1101;
	mem[1093] = 4'b1110;
	mem[1094] = 4'b0111;
	mem[1095] = 4'b0010;
	mem[1096] = 4'b0001;
	mem[1097] = 4'b0001;
	mem[1098] = 4'b0010;
	mem[1099] = 4'b0010;
	mem[1100] = 4'b0010;
	mem[1101] = 4'b0010;
	mem[1102] = 4'b0010;
	mem[1103] = 4'b0011;
	mem[1104] = 4'b0011;
	mem[1105] = 4'b0010;
	mem[1106] = 4'b0010;
	mem[1107] = 4'b0010;
	mem[1108] = 4'b0010;
	mem[1109] = 4'b0011;
	mem[1110] = 4'b0011;
	mem[1111] = 4'b0011;
	mem[1112] = 4'b0011;
	mem[1113] = 4'b0011;
	mem[1114] = 4'b0011;
	mem[1115] = 4'b0011;
	mem[1116] = 4'b0011;
	mem[1117] = 4'b0011;
	mem[1118] = 4'b0100;
	mem[1119] = 4'b0100;
	mem[1120] = 4'b0100;
	mem[1121] = 4'b0100;
	mem[1122] = 4'b0100;
	mem[1123] = 4'b0100;
	mem[1124] = 4'b0100;
	mem[1125] = 4'b0100;
	mem[1126] = 4'b0100;
	mem[1127] = 4'b0101;
	mem[1128] = 4'b0101;
	mem[1129] = 4'b0101;
	mem[1130] = 4'b0101;
	mem[1131] = 4'b0101;
	mem[1132] = 4'b0101;
	mem[1133] = 4'b0101;
	mem[1134] = 4'b0101;
	mem[1135] = 4'b0101;
	mem[1136] = 4'b0101;
	mem[1137] = 4'b0110;
	mem[1138] = 4'b0110;
	mem[1139] = 4'b0110;
	mem[1140] = 4'b0110;
	mem[1141] = 4'b0110;
	mem[1142] = 4'b0110;
	mem[1143] = 4'b0110;
	mem[1144] = 4'b0110;
	mem[1145] = 4'b0110;
	mem[1146] = 4'b0001;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0000;
	mem[1156] = 4'b0000;
	mem[1157] = 4'b0000;
	mem[1158] = 4'b0000;
	mem[1159] = 4'b0000;
	mem[1160] = 4'b0000;
	mem[1161] = 4'b0001;
	mem[1162] = 4'b0001;
	mem[1163] = 4'b0001;
	mem[1164] = 4'b0001;
	mem[1165] = 4'b0001;
	mem[1166] = 4'b0010;
	mem[1167] = 4'b0011;
	mem[1168] = 4'b0011;
	mem[1169] = 4'b0011;
	mem[1170] = 4'b0100;
	mem[1171] = 4'b0011;
	mem[1172] = 4'b0100;
	mem[1173] = 4'b0101;
	mem[1174] = 4'b0101;
	mem[1175] = 4'b0100;
	mem[1176] = 4'b0100;
	mem[1177] = 4'b0101;
	mem[1178] = 4'b0110;
	mem[1179] = 4'b0110;
	mem[1180] = 4'b0110;
	mem[1181] = 4'b0110;
	mem[1182] = 4'b0110;
	mem[1183] = 4'b0111;
	mem[1184] = 4'b1000;
	mem[1185] = 4'b1000;
	mem[1186] = 4'b1000;
	mem[1187] = 4'b1000;
	mem[1188] = 4'b1000;
	mem[1189] = 4'b1001;
	mem[1190] = 4'b1001;
	mem[1191] = 4'b1001;
	mem[1192] = 4'b1001;
	mem[1193] = 4'b1001;
	mem[1194] = 4'b1010;
	mem[1195] = 4'b1011;
	mem[1196] = 4'b1011;
	mem[1197] = 4'b1011;
	mem[1198] = 4'b1011;
	mem[1199] = 4'b1011;
	mem[1200] = 4'b1100;
	mem[1201] = 4'b1100;
	mem[1202] = 4'b1100;
	mem[1203] = 4'b1100;
	mem[1204] = 4'b1100;
	mem[1205] = 4'b1101;
	mem[1206] = 4'b1110;
	mem[1207] = 4'b1110;
	mem[1208] = 4'b1110;
	mem[1209] = 4'b1110;
	mem[1210] = 4'b1110;
	mem[1211] = 4'b1111;
	mem[1212] = 4'b1111;
	mem[1213] = 4'b1111;
	mem[1214] = 4'b1111;
	mem[1215] = 4'b1111;
	mem[1216] = 4'b1111;
	mem[1217] = 4'b1111;
	mem[1218] = 4'b1111;
	mem[1219] = 4'b1101;
	mem[1220] = 4'b1110;
	mem[1221] = 4'b1111;
	mem[1222] = 4'b0111;
	mem[1223] = 4'b0001;
	mem[1224] = 4'b0010;
	mem[1225] = 4'b0010;
	mem[1226] = 4'b0010;
	mem[1227] = 4'b0011;
	mem[1228] = 4'b0010;
	mem[1229] = 4'b0010;
	mem[1230] = 4'b0011;
	mem[1231] = 4'b0011;
	mem[1232] = 4'b0011;
	mem[1233] = 4'b0010;
	mem[1234] = 4'b0010;
	mem[1235] = 4'b0011;
	mem[1236] = 4'b0011;
	mem[1237] = 4'b0011;
	mem[1238] = 4'b0011;
	mem[1239] = 4'b0011;
	mem[1240] = 4'b0011;
	mem[1241] = 4'b0011;
	mem[1242] = 4'b0011;
	mem[1243] = 4'b0011;
	mem[1244] = 4'b0100;
	mem[1245] = 4'b0100;
	mem[1246] = 4'b0100;
	mem[1247] = 4'b0100;
	mem[1248] = 4'b0100;
	mem[1249] = 4'b0100;
	mem[1250] = 4'b0100;
	mem[1251] = 4'b0100;
	mem[1252] = 4'b0100;
	mem[1253] = 4'b0101;
	mem[1254] = 4'b0101;
	mem[1255] = 4'b0101;
	mem[1256] = 4'b0101;
	mem[1257] = 4'b0101;
	mem[1258] = 4'b0101;
	mem[1259] = 4'b0101;
	mem[1260] = 4'b0101;
	mem[1261] = 4'b0101;
	mem[1262] = 4'b0110;
	mem[1263] = 4'b0110;
	mem[1264] = 4'b0110;
	mem[1265] = 4'b0110;
	mem[1266] = 4'b0110;
	mem[1267] = 4'b0110;
	mem[1268] = 4'b0110;
	mem[1269] = 4'b0110;
	mem[1270] = 4'b0110;
	mem[1271] = 4'b0111;
	mem[1272] = 4'b0111;
	mem[1273] = 4'b0110;
	mem[1274] = 4'b0001;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0000;
	mem[1284] = 4'b0000;
	mem[1285] = 4'b0000;
	mem[1286] = 4'b0000;
	mem[1287] = 4'b0000;
	mem[1288] = 4'b0000;
	mem[1289] = 4'b0001;
	mem[1290] = 4'b0001;
	mem[1291] = 4'b0001;
	mem[1292] = 4'b0001;
	mem[1293] = 4'b0001;
	mem[1294] = 4'b0010;
	mem[1295] = 4'b0011;
	mem[1296] = 4'b0011;
	mem[1297] = 4'b0100;
	mem[1298] = 4'b0011;
	mem[1299] = 4'b0011;
	mem[1300] = 4'b0100;
	mem[1301] = 4'b0100;
	mem[1302] = 4'b0100;
	mem[1303] = 4'b0100;
	mem[1304] = 4'b0100;
	mem[1305] = 4'b0101;
	mem[1306] = 4'b0110;
	mem[1307] = 4'b0101;
	mem[1308] = 4'b0110;
	mem[1309] = 4'b0110;
	mem[1310] = 4'b0110;
	mem[1311] = 4'b0111;
	mem[1312] = 4'b1000;
	mem[1313] = 4'b1000;
	mem[1314] = 4'b1000;
	mem[1315] = 4'b1000;
	mem[1316] = 4'b1000;
	mem[1317] = 4'b1001;
	mem[1318] = 4'b1001;
	mem[1319] = 4'b1001;
	mem[1320] = 4'b1001;
	mem[1321] = 4'b1001;
	mem[1322] = 4'b1010;
	mem[1323] = 4'b1011;
	mem[1324] = 4'b1011;
	mem[1325] = 4'b1011;
	mem[1326] = 4'b1011;
	mem[1327] = 4'b1011;
	mem[1328] = 4'b1100;
	mem[1329] = 4'b1100;
	mem[1330] = 4'b1100;
	mem[1331] = 4'b1100;
	mem[1332] = 4'b1100;
	mem[1333] = 4'b1101;
	mem[1334] = 4'b1110;
	mem[1335] = 4'b1110;
	mem[1336] = 4'b1110;
	mem[1337] = 4'b1110;
	mem[1338] = 4'b1110;
	mem[1339] = 4'b1111;
	mem[1340] = 4'b1111;
	mem[1341] = 4'b1111;
	mem[1342] = 4'b1111;
	mem[1343] = 4'b1111;
	mem[1344] = 4'b1111;
	mem[1345] = 4'b1111;
	mem[1346] = 4'b1110;
	mem[1347] = 4'b1101;
	mem[1348] = 4'b1110;
	mem[1349] = 4'b1111;
	mem[1350] = 4'b0111;
	mem[1351] = 4'b0010;
	mem[1352] = 4'b0010;
	mem[1353] = 4'b0010;
	mem[1354] = 4'b0010;
	mem[1355] = 4'b0011;
	mem[1356] = 4'b0011;
	mem[1357] = 4'b0010;
	mem[1358] = 4'b0010;
	mem[1359] = 4'b0011;
	mem[1360] = 4'b0011;
	mem[1361] = 4'b0011;
	mem[1362] = 4'b0011;
	mem[1363] = 4'b0011;
	mem[1364] = 4'b0011;
	mem[1365] = 4'b0011;
	mem[1366] = 4'b0011;
	mem[1367] = 4'b0011;
	mem[1368] = 4'b0011;
	mem[1369] = 4'b0100;
	mem[1370] = 4'b0100;
	mem[1371] = 4'b0100;
	mem[1372] = 4'b0100;
	mem[1373] = 4'b0100;
	mem[1374] = 4'b0100;
	mem[1375] = 4'b0100;
	mem[1376] = 4'b0100;
	mem[1377] = 4'b0100;
	mem[1378] = 4'b0101;
	mem[1379] = 4'b0101;
	mem[1380] = 4'b0101;
	mem[1381] = 4'b0101;
	mem[1382] = 4'b0101;
	mem[1383] = 4'b0101;
	mem[1384] = 4'b0101;
	mem[1385] = 4'b0101;
	mem[1386] = 4'b0101;
	mem[1387] = 4'b0110;
	mem[1388] = 4'b0110;
	mem[1389] = 4'b0110;
	mem[1390] = 4'b0110;
	mem[1391] = 4'b0110;
	mem[1392] = 4'b0110;
	mem[1393] = 4'b0110;
	mem[1394] = 4'b0110;
	mem[1395] = 4'b0110;
	mem[1396] = 4'b0110;
	mem[1397] = 4'b0111;
	mem[1398] = 4'b0111;
	mem[1399] = 4'b0111;
	mem[1400] = 4'b0111;
	mem[1401] = 4'b0111;
	mem[1402] = 4'b0001;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0000;
	mem[1412] = 4'b0000;
	mem[1413] = 4'b0000;
	mem[1414] = 4'b0000;
	mem[1415] = 4'b0000;
	mem[1416] = 4'b0000;
	mem[1417] = 4'b0001;
	mem[1418] = 4'b0001;
	mem[1419] = 4'b0001;
	mem[1420] = 4'b0001;
	mem[1421] = 4'b0001;
	mem[1422] = 4'b0010;
	mem[1423] = 4'b0011;
	mem[1424] = 4'b0011;
	mem[1425] = 4'b0100;
	mem[1426] = 4'b0011;
	mem[1427] = 4'b0011;
	mem[1428] = 4'b0100;
	mem[1429] = 4'b0100;
	mem[1430] = 4'b0100;
	mem[1431] = 4'b0100;
	mem[1432] = 4'b0100;
	mem[1433] = 4'b0101;
	mem[1434] = 4'b0101;
	mem[1435] = 4'b0101;
	mem[1436] = 4'b0110;
	mem[1437] = 4'b0110;
	mem[1438] = 4'b0110;
	mem[1439] = 4'b0111;
	mem[1440] = 4'b1000;
	mem[1441] = 4'b1000;
	mem[1442] = 4'b1000;
	mem[1443] = 4'b1000;
	mem[1444] = 4'b1000;
	mem[1445] = 4'b1001;
	mem[1446] = 4'b1001;
	mem[1447] = 4'b1001;
	mem[1448] = 4'b1001;
	mem[1449] = 4'b1001;
	mem[1450] = 4'b1010;
	mem[1451] = 4'b1011;
	mem[1452] = 4'b1011;
	mem[1453] = 4'b1011;
	mem[1454] = 4'b1011;
	mem[1455] = 4'b1011;
	mem[1456] = 4'b1100;
	mem[1457] = 4'b1100;
	mem[1458] = 4'b1100;
	mem[1459] = 4'b1100;
	mem[1460] = 4'b1100;
	mem[1461] = 4'b1101;
	mem[1462] = 4'b1110;
	mem[1463] = 4'b1110;
	mem[1464] = 4'b1110;
	mem[1465] = 4'b1110;
	mem[1466] = 4'b1110;
	mem[1467] = 4'b1111;
	mem[1468] = 4'b1111;
	mem[1469] = 4'b1111;
	mem[1470] = 4'b1111;
	mem[1471] = 4'b1111;
	mem[1472] = 4'b1111;
	mem[1473] = 4'b1111;
	mem[1474] = 4'b1110;
	mem[1475] = 4'b1101;
	mem[1476] = 4'b1110;
	mem[1477] = 4'b1111;
	mem[1478] = 4'b0111;
	mem[1479] = 4'b0010;
	mem[1480] = 4'b0010;
	mem[1481] = 4'b0010;
	mem[1482] = 4'b0010;
	mem[1483] = 4'b0011;
	mem[1484] = 4'b0011;
	mem[1485] = 4'b0011;
	mem[1486] = 4'b0011;
	mem[1487] = 4'b0011;
	mem[1488] = 4'b0011;
	mem[1489] = 4'b0011;
	mem[1490] = 4'b0011;
	mem[1491] = 4'b0011;
	mem[1492] = 4'b0011;
	mem[1493] = 4'b0011;
	mem[1494] = 4'b0011;
	mem[1495] = 4'b0100;
	mem[1496] = 4'b0100;
	mem[1497] = 4'b0100;
	mem[1498] = 4'b0100;
	mem[1499] = 4'b0100;
	mem[1500] = 4'b0100;
	mem[1501] = 4'b0100;
	mem[1502] = 4'b0100;
	mem[1503] = 4'b0100;
	mem[1504] = 4'b0101;
	mem[1505] = 4'b0101;
	mem[1506] = 4'b0101;
	mem[1507] = 4'b0101;
	mem[1508] = 4'b0101;
	mem[1509] = 4'b0101;
	mem[1510] = 4'b0101;
	mem[1511] = 4'b0101;
	mem[1512] = 4'b0101;
	mem[1513] = 4'b0110;
	mem[1514] = 4'b0110;
	mem[1515] = 4'b0110;
	mem[1516] = 4'b0110;
	mem[1517] = 4'b0110;
	mem[1518] = 4'b0110;
	mem[1519] = 4'b0110;
	mem[1520] = 4'b0110;
	mem[1521] = 4'b0110;
	mem[1522] = 4'b0111;
	mem[1523] = 4'b0111;
	mem[1524] = 4'b0111;
	mem[1525] = 4'b0111;
	mem[1526] = 4'b0111;
	mem[1527] = 4'b0111;
	mem[1528] = 4'b0111;
	mem[1529] = 4'b0111;
	mem[1530] = 4'b0001;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0000;
	mem[1540] = 4'b0000;
	mem[1541] = 4'b0000;
	mem[1542] = 4'b0000;
	mem[1543] = 4'b0000;
	mem[1544] = 4'b0000;
	mem[1545] = 4'b0001;
	mem[1546] = 4'b0001;
	mem[1547] = 4'b0001;
	mem[1548] = 4'b0001;
	mem[1549] = 4'b0001;
	mem[1550] = 4'b0010;
	mem[1551] = 4'b0010;
	mem[1552] = 4'b0010;
	mem[1553] = 4'b0011;
	mem[1554] = 4'b0010;
	mem[1555] = 4'b0010;
	mem[1556] = 4'b0100;
	mem[1557] = 4'b0100;
	mem[1558] = 4'b0100;
	mem[1559] = 4'b0100;
	mem[1560] = 4'b0100;
	mem[1561] = 4'b0100;
	mem[1562] = 4'b0101;
	mem[1563] = 4'b0101;
	mem[1564] = 4'b0101;
	mem[1565] = 4'b0110;
	mem[1566] = 4'b0101;
	mem[1567] = 4'b0110;
	mem[1568] = 4'b0111;
	mem[1569] = 4'b0111;
	mem[1570] = 4'b0111;
	mem[1571] = 4'b0111;
	mem[1572] = 4'b0111;
	mem[1573] = 4'b1000;
	mem[1574] = 4'b1000;
	mem[1575] = 4'b1000;
	mem[1576] = 4'b1000;
	mem[1577] = 4'b1000;
	mem[1578] = 4'b1001;
	mem[1579] = 4'b1010;
	mem[1580] = 4'b1010;
	mem[1581] = 4'b1010;
	mem[1582] = 4'b1010;
	mem[1583] = 4'b1010;
	mem[1584] = 4'b1011;
	mem[1585] = 4'b1011;
	mem[1586] = 4'b1011;
	mem[1587] = 4'b1011;
	mem[1588] = 4'b1011;
	mem[1589] = 4'b1100;
	mem[1590] = 4'b1101;
	mem[1591] = 4'b1101;
	mem[1592] = 4'b1101;
	mem[1593] = 4'b1101;
	mem[1594] = 4'b1101;
	mem[1595] = 4'b1101;
	mem[1596] = 4'b1101;
	mem[1597] = 4'b1101;
	mem[1598] = 4'b1101;
	mem[1599] = 4'b1101;
	mem[1600] = 4'b1101;
	mem[1601] = 4'b1110;
	mem[1602] = 4'b1110;
	mem[1603] = 4'b1100;
	mem[1604] = 4'b1100;
	mem[1605] = 4'b1101;
	mem[1606] = 4'b0111;
	mem[1607] = 4'b0010;
	mem[1608] = 4'b0010;
	mem[1609] = 4'b0010;
	mem[1610] = 4'b0010;
	mem[1611] = 4'b0011;
	mem[1612] = 4'b0011;
	mem[1613] = 4'b0010;
	mem[1614] = 4'b0011;
	mem[1615] = 4'b0011;
	mem[1616] = 4'b0011;
	mem[1617] = 4'b0011;
	mem[1618] = 4'b0011;
	mem[1619] = 4'b0011;
	mem[1620] = 4'b0011;
	mem[1621] = 4'b0011;
	mem[1622] = 4'b0011;
	mem[1623] = 4'b0011;
	mem[1624] = 4'b0100;
	mem[1625] = 4'b0100;
	mem[1626] = 4'b0100;
	mem[1627] = 4'b0100;
	mem[1628] = 4'b0100;
	mem[1629] = 4'b0100;
	mem[1630] = 4'b0100;
	mem[1631] = 4'b0100;
	mem[1632] = 4'b0100;
	mem[1633] = 4'b0100;
	mem[1634] = 4'b0101;
	mem[1635] = 4'b0101;
	mem[1636] = 4'b0101;
	mem[1637] = 4'b0101;
	mem[1638] = 4'b0101;
	mem[1639] = 4'b0101;
	mem[1640] = 4'b0101;
	mem[1641] = 4'b0101;
	mem[1642] = 4'b0101;
	mem[1643] = 4'b0101;
	mem[1644] = 4'b0110;
	mem[1645] = 4'b0110;
	mem[1646] = 4'b0110;
	mem[1647] = 4'b0110;
	mem[1648] = 4'b0110;
	mem[1649] = 4'b0110;
	mem[1650] = 4'b0110;
	mem[1651] = 4'b0110;
	mem[1652] = 4'b0110;
	mem[1653] = 4'b0110;
	mem[1654] = 4'b0111;
	mem[1655] = 4'b0111;
	mem[1656] = 4'b0111;
	mem[1657] = 4'b0111;
	mem[1658] = 4'b0001;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0000;
	mem[1668] = 4'b0000;
	mem[1669] = 4'b0000;
	mem[1670] = 4'b0000;
	mem[1671] = 4'b0000;
	mem[1672] = 4'b0000;
	mem[1673] = 4'b0000;
	mem[1674] = 4'b0000;
	mem[1675] = 4'b0000;
	mem[1676] = 4'b0000;
	mem[1677] = 4'b0000;
	mem[1678] = 4'b0000;
	mem[1679] = 4'b0000;
	mem[1680] = 4'b0000;
	mem[1681] = 4'b0001;
	mem[1682] = 4'b0000;
	mem[1683] = 4'b0000;
	mem[1684] = 4'b0000;
	mem[1685] = 4'b0000;
	mem[1686] = 4'b0000;
	mem[1687] = 4'b0000;
	mem[1688] = 4'b0000;
	mem[1689] = 4'b0001;
	mem[1690] = 4'b0000;
	mem[1691] = 4'b0001;
	mem[1692] = 4'b0001;
	mem[1693] = 4'b0001;
	mem[1694] = 4'b0000;
	mem[1695] = 4'b0000;
	mem[1696] = 4'b0000;
	mem[1697] = 4'b0000;
	mem[1698] = 4'b0000;
	mem[1699] = 4'b0000;
	mem[1700] = 4'b0000;
	mem[1701] = 4'b0000;
	mem[1702] = 4'b0000;
	mem[1703] = 4'b0000;
	mem[1704] = 4'b0000;
	mem[1705] = 4'b0000;
	mem[1706] = 4'b0000;
	mem[1707] = 4'b0001;
	mem[1708] = 4'b0001;
	mem[1709] = 4'b0001;
	mem[1710] = 4'b0001;
	mem[1711] = 4'b0001;
	mem[1712] = 4'b0001;
	mem[1713] = 4'b0001;
	mem[1714] = 4'b0001;
	mem[1715] = 4'b0001;
	mem[1716] = 4'b0001;
	mem[1717] = 4'b0001;
	mem[1718] = 4'b0001;
	mem[1719] = 4'b0001;
	mem[1720] = 4'b0001;
	mem[1721] = 4'b0001;
	mem[1722] = 4'b0001;
	mem[1723] = 4'b0001;
	mem[1724] = 4'b0001;
	mem[1725] = 4'b0001;
	mem[1726] = 4'b0001;
	mem[1727] = 4'b0001;
	mem[1728] = 4'b0001;
	mem[1729] = 4'b0010;
	mem[1730] = 4'b0001;
	mem[1731] = 4'b0010;
	mem[1732] = 4'b0001;
	mem[1733] = 4'b0001;
	mem[1734] = 4'b0001;
	mem[1735] = 4'b0000;
	mem[1736] = 4'b0000;
	mem[1737] = 4'b0000;
	mem[1738] = 4'b0001;
	mem[1739] = 4'b0001;
	mem[1740] = 4'b0000;
	mem[1741] = 4'b0000;
	mem[1742] = 4'b0000;
	mem[1743] = 4'b0000;
	mem[1744] = 4'b0000;
	mem[1745] = 4'b0000;
	mem[1746] = 4'b0000;
	mem[1747] = 4'b0000;
	mem[1748] = 4'b0000;
	mem[1749] = 4'b0000;
	mem[1750] = 4'b0000;
	mem[1751] = 4'b0000;
	mem[1752] = 4'b0000;
	mem[1753] = 4'b0000;
	mem[1754] = 4'b0000;
	mem[1755] = 4'b0000;
	mem[1756] = 4'b0000;
	mem[1757] = 4'b0000;
	mem[1758] = 4'b0000;
	mem[1759] = 4'b0000;
	mem[1760] = 4'b0000;
	mem[1761] = 4'b0000;
	mem[1762] = 4'b0000;
	mem[1763] = 4'b0000;
	mem[1764] = 4'b0000;
	mem[1765] = 4'b0000;
	mem[1766] = 4'b0000;
	mem[1767] = 4'b0000;
	mem[1768] = 4'b0000;
	mem[1769] = 4'b0000;
	mem[1770] = 4'b0000;
	mem[1771] = 4'b0000;
	mem[1772] = 4'b0000;
	mem[1773] = 4'b0000;
	mem[1774] = 4'b0000;
	mem[1775] = 4'b0000;
	mem[1776] = 4'b0000;
	mem[1777] = 4'b0000;
	mem[1778] = 4'b0000;
	mem[1779] = 4'b0000;
	mem[1780] = 4'b0000;
	mem[1781] = 4'b0000;
	mem[1782] = 4'b0000;
	mem[1783] = 4'b0000;
	mem[1784] = 4'b0000;
	mem[1785] = 4'b0000;
	mem[1786] = 4'b0000;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0000;
	mem[1796] = 4'b0000;
	mem[1797] = 4'b0000;
	mem[1798] = 4'b0000;
	mem[1799] = 4'b0000;
	mem[1800] = 4'b0000;
	mem[1801] = 4'b0000;
	mem[1802] = 4'b0000;
	mem[1803] = 4'b0000;
	mem[1804] = 4'b0000;
	mem[1805] = 4'b0000;
	mem[1806] = 4'b0000;
	mem[1807] = 4'b0000;
	mem[1808] = 4'b0000;
	mem[1809] = 4'b0000;
	mem[1810] = 4'b0001;
	mem[1811] = 4'b0000;
	mem[1812] = 4'b0000;
	mem[1813] = 4'b0000;
	mem[1814] = 4'b0000;
	mem[1815] = 4'b0000;
	mem[1816] = 4'b0000;
	mem[1817] = 4'b0000;
	mem[1818] = 4'b0000;
	mem[1819] = 4'b0000;
	mem[1820] = 4'b0000;
	mem[1821] = 4'b0001;
	mem[1822] = 4'b0000;
	mem[1823] = 4'b0000;
	mem[1824] = 4'b0000;
	mem[1825] = 4'b0000;
	mem[1826] = 4'b0000;
	mem[1827] = 4'b0000;
	mem[1828] = 4'b0000;
	mem[1829] = 4'b0000;
	mem[1830] = 4'b0000;
	mem[1831] = 4'b0000;
	mem[1832] = 4'b0000;
	mem[1833] = 4'b0000;
	mem[1834] = 4'b0000;
	mem[1835] = 4'b0000;
	mem[1836] = 4'b0000;
	mem[1837] = 4'b0000;
	mem[1838] = 4'b0000;
	mem[1839] = 4'b0000;
	mem[1840] = 4'b0000;
	mem[1841] = 4'b0000;
	mem[1842] = 4'b0000;
	mem[1843] = 4'b0000;
	mem[1844] = 4'b0000;
	mem[1845] = 4'b0000;
	mem[1846] = 4'b0000;
	mem[1847] = 4'b0000;
	mem[1848] = 4'b0000;
	mem[1849] = 4'b0000;
	mem[1850] = 4'b0000;
	mem[1851] = 4'b0000;
	mem[1852] = 4'b0000;
	mem[1853] = 4'b0000;
	mem[1854] = 4'b0000;
	mem[1855] = 4'b0000;
	mem[1856] = 4'b0000;
	mem[1857] = 4'b0001;
	mem[1858] = 4'b0000;
	mem[1859] = 4'b0000;
	mem[1860] = 4'b0000;
	mem[1861] = 4'b0000;
	mem[1862] = 4'b0000;
	mem[1863] = 4'b0000;
	mem[1864] = 4'b0000;
	mem[1865] = 4'b0001;
	mem[1866] = 4'b0001;
	mem[1867] = 4'b0000;
	mem[1868] = 4'b0000;
	mem[1869] = 4'b0000;
	mem[1870] = 4'b0000;
	mem[1871] = 4'b0000;
	mem[1872] = 4'b0000;
	mem[1873] = 4'b0000;
	mem[1874] = 4'b0000;
	mem[1875] = 4'b0000;
	mem[1876] = 4'b0000;
	mem[1877] = 4'b0000;
	mem[1878] = 4'b0000;
	mem[1879] = 4'b0000;
	mem[1880] = 4'b0000;
	mem[1881] = 4'b0000;
	mem[1882] = 4'b0000;
	mem[1883] = 4'b0000;
	mem[1884] = 4'b0000;
	mem[1885] = 4'b0000;
	mem[1886] = 4'b0000;
	mem[1887] = 4'b0000;
	mem[1888] = 4'b0000;
	mem[1889] = 4'b0000;
	mem[1890] = 4'b0000;
	mem[1891] = 4'b0000;
	mem[1892] = 4'b0000;
	mem[1893] = 4'b0000;
	mem[1894] = 4'b0000;
	mem[1895] = 4'b0000;
	mem[1896] = 4'b0000;
	mem[1897] = 4'b0000;
	mem[1898] = 4'b0000;
	mem[1899] = 4'b0000;
	mem[1900] = 4'b0000;
	mem[1901] = 4'b0000;
	mem[1902] = 4'b0000;
	mem[1903] = 4'b0000;
	mem[1904] = 4'b0000;
	mem[1905] = 4'b0000;
	mem[1906] = 4'b0000;
	mem[1907] = 4'b0000;
	mem[1908] = 4'b0000;
	mem[1909] = 4'b0000;
	mem[1910] = 4'b0000;
	mem[1911] = 4'b0000;
	mem[1912] = 4'b0000;
	mem[1913] = 4'b0000;
	mem[1914] = 4'b0000;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0000;
	mem[1924] = 4'b0000;
	mem[1925] = 4'b0000;
	mem[1926] = 4'b0000;
	mem[1927] = 4'b0000;
	mem[1928] = 4'b0000;
	mem[1929] = 4'b0000;
	mem[1930] = 4'b0000;
	mem[1931] = 4'b0000;
	mem[1932] = 4'b0000;
	mem[1933] = 4'b0000;
	mem[1934] = 4'b0000;
	mem[1935] = 4'b0000;
	mem[1936] = 4'b0000;
	mem[1937] = 4'b0000;
	mem[1938] = 4'b0000;
	mem[1939] = 4'b0000;
	mem[1940] = 4'b0000;
	mem[1941] = 4'b0000;
	mem[1942] = 4'b0000;
	mem[1943] = 4'b0000;
	mem[1944] = 4'b0000;
	mem[1945] = 4'b0000;
	mem[1946] = 4'b0000;
	mem[1947] = 4'b0000;
	mem[1948] = 4'b0001;
	mem[1949] = 4'b0000;
	mem[1950] = 4'b0000;
	mem[1951] = 4'b0000;
	mem[1952] = 4'b0000;
	mem[1953] = 4'b0000;
	mem[1954] = 4'b0000;
	mem[1955] = 4'b0000;
	mem[1956] = 4'b0000;
	mem[1957] = 4'b0000;
	mem[1958] = 4'b0000;
	mem[1959] = 4'b0000;
	mem[1960] = 4'b0000;
	mem[1961] = 4'b0000;
	mem[1962] = 4'b0000;
	mem[1963] = 4'b0000;
	mem[1964] = 4'b0000;
	mem[1965] = 4'b0000;
	mem[1966] = 4'b0000;
	mem[1967] = 4'b0000;
	mem[1968] = 4'b0000;
	mem[1969] = 4'b0000;
	mem[1970] = 4'b0000;
	mem[1971] = 4'b0000;
	mem[1972] = 4'b0000;
	mem[1973] = 4'b0000;
	mem[1974] = 4'b0000;
	mem[1975] = 4'b0000;
	mem[1976] = 4'b0000;
	mem[1977] = 4'b0000;
	mem[1978] = 4'b0000;
	mem[1979] = 4'b0000;
	mem[1980] = 4'b0000;
	mem[1981] = 4'b0000;
	mem[1982] = 4'b0001;
	mem[1983] = 4'b0001;
	mem[1984] = 4'b0001;
	mem[1985] = 4'b0000;
	mem[1986] = 4'b0000;
	mem[1987] = 4'b0000;
	mem[1988] = 4'b0000;
	mem[1989] = 4'b0000;
	mem[1990] = 4'b0001;
	mem[1991] = 4'b0001;
	mem[1992] = 4'b0001;
	mem[1993] = 4'b0001;
	mem[1994] = 4'b0000;
	mem[1995] = 4'b0000;
	mem[1996] = 4'b0000;
	mem[1997] = 4'b0000;
	mem[1998] = 4'b0000;
	mem[1999] = 4'b0000;
	mem[2000] = 4'b0000;
	mem[2001] = 4'b0000;
	mem[2002] = 4'b0000;
	mem[2003] = 4'b0000;
	mem[2004] = 4'b0000;
	mem[2005] = 4'b0000;
	mem[2006] = 4'b0000;
	mem[2007] = 4'b0000;
	mem[2008] = 4'b0000;
	mem[2009] = 4'b0000;
	mem[2010] = 4'b0000;
	mem[2011] = 4'b0000;
	mem[2012] = 4'b0000;
	mem[2013] = 4'b0000;
	mem[2014] = 4'b0000;
	mem[2015] = 4'b0000;
	mem[2016] = 4'b0000;
	mem[2017] = 4'b0000;
	mem[2018] = 4'b0000;
	mem[2019] = 4'b0000;
	mem[2020] = 4'b0000;
	mem[2021] = 4'b0000;
	mem[2022] = 4'b0000;
	mem[2023] = 4'b0000;
	mem[2024] = 4'b0000;
	mem[2025] = 4'b0000;
	mem[2026] = 4'b0000;
	mem[2027] = 4'b0000;
	mem[2028] = 4'b0000;
	mem[2029] = 4'b0000;
	mem[2030] = 4'b0000;
	mem[2031] = 4'b0000;
	mem[2032] = 4'b0000;
	mem[2033] = 4'b0000;
	mem[2034] = 4'b0000;
	mem[2035] = 4'b0000;
	mem[2036] = 4'b0000;
	mem[2037] = 4'b0000;
	mem[2038] = 4'b0000;
	mem[2039] = 4'b0000;
	mem[2040] = 4'b0000;
	mem[2041] = 4'b0000;
	mem[2042] = 4'b0000;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0000;
	mem[2052] = 4'b0000;
	mem[2053] = 4'b0000;
	mem[2054] = 4'b0000;
	mem[2055] = 4'b0000;
	mem[2056] = 4'b0000;
	mem[2057] = 4'b0000;
	mem[2058] = 4'b0000;
	mem[2059] = 4'b0000;
	mem[2060] = 4'b0000;
	mem[2061] = 4'b0000;
	mem[2062] = 4'b0000;
	mem[2063] = 4'b0000;
	mem[2064] = 4'b0000;
	mem[2065] = 4'b0000;
	mem[2066] = 4'b0000;
	mem[2067] = 4'b0000;
	mem[2068] = 4'b0000;
	mem[2069] = 4'b0000;
	mem[2070] = 4'b0000;
	mem[2071] = 4'b0000;
	mem[2072] = 4'b0000;
	mem[2073] = 4'b0000;
	mem[2074] = 4'b0000;
	mem[2075] = 4'b0000;
	mem[2076] = 4'b0001;
	mem[2077] = 4'b0000;
	mem[2078] = 4'b0000;
	mem[2079] = 4'b0000;
	mem[2080] = 4'b0000;
	mem[2081] = 4'b0000;
	mem[2082] = 4'b0000;
	mem[2083] = 4'b0000;
	mem[2084] = 4'b0000;
	mem[2085] = 4'b0000;
	mem[2086] = 4'b0000;
	mem[2087] = 4'b0000;
	mem[2088] = 4'b0000;
	mem[2089] = 4'b0000;
	mem[2090] = 4'b0000;
	mem[2091] = 4'b0000;
	mem[2092] = 4'b0000;
	mem[2093] = 4'b0000;
	mem[2094] = 4'b0000;
	mem[2095] = 4'b0000;
	mem[2096] = 4'b0000;
	mem[2097] = 4'b0000;
	mem[2098] = 4'b0000;
	mem[2099] = 4'b0000;
	mem[2100] = 4'b0000;
	mem[2101] = 4'b0000;
	mem[2102] = 4'b0000;
	mem[2103] = 4'b0000;
	mem[2104] = 4'b0000;
	mem[2105] = 4'b0000;
	mem[2106] = 4'b0000;
	mem[2107] = 4'b0000;
	mem[2108] = 4'b0000;
	mem[2109] = 4'b0000;
	mem[2110] = 4'b0001;
	mem[2111] = 4'b0000;
	mem[2112] = 4'b0000;
	mem[2113] = 4'b0000;
	mem[2114] = 4'b0000;
	mem[2115] = 4'b0000;
	mem[2116] = 4'b0000;
	mem[2117] = 4'b0000;
	mem[2118] = 4'b0000;
	mem[2119] = 4'b0000;
	mem[2120] = 4'b0000;
	mem[2121] = 4'b0000;
	mem[2122] = 4'b0000;
	mem[2123] = 4'b0000;
	mem[2124] = 4'b0000;
	mem[2125] = 4'b0000;
	mem[2126] = 4'b0000;
	mem[2127] = 4'b0000;
	mem[2128] = 4'b0000;
	mem[2129] = 4'b0000;
	mem[2130] = 4'b0000;
	mem[2131] = 4'b0000;
	mem[2132] = 4'b0000;
	mem[2133] = 4'b0000;
	mem[2134] = 4'b0000;
	mem[2135] = 4'b0000;
	mem[2136] = 4'b0000;
	mem[2137] = 4'b0000;
	mem[2138] = 4'b0000;
	mem[2139] = 4'b0000;
	mem[2140] = 4'b0000;
	mem[2141] = 4'b0000;
	mem[2142] = 4'b0000;
	mem[2143] = 4'b0000;
	mem[2144] = 4'b0000;
	mem[2145] = 4'b0000;
	mem[2146] = 4'b0000;
	mem[2147] = 4'b0000;
	mem[2148] = 4'b0000;
	mem[2149] = 4'b0000;
	mem[2150] = 4'b0000;
	mem[2151] = 4'b0000;
	mem[2152] = 4'b0000;
	mem[2153] = 4'b0000;
	mem[2154] = 4'b0000;
	mem[2155] = 4'b0000;
	mem[2156] = 4'b0000;
	mem[2157] = 4'b0000;
	mem[2158] = 4'b0000;
	mem[2159] = 4'b0000;
	mem[2160] = 4'b0000;
	mem[2161] = 4'b0000;
	mem[2162] = 4'b0000;
	mem[2163] = 4'b0000;
	mem[2164] = 4'b0000;
	mem[2165] = 4'b0000;
	mem[2166] = 4'b0000;
	mem[2167] = 4'b0000;
	mem[2168] = 4'b0000;
	mem[2169] = 4'b0000;
	mem[2170] = 4'b0000;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0000;
	mem[2180] = 4'b0000;
	mem[2181] = 4'b0000;
	mem[2182] = 4'b0000;
	mem[2183] = 4'b0000;
	mem[2184] = 4'b0000;
	mem[2185] = 4'b0000;
	mem[2186] = 4'b0000;
	mem[2187] = 4'b0000;
	mem[2188] = 4'b0000;
	mem[2189] = 4'b0000;
	mem[2190] = 4'b0000;
	mem[2191] = 4'b0000;
	mem[2192] = 4'b0000;
	mem[2193] = 4'b0000;
	mem[2194] = 4'b0000;
	mem[2195] = 4'b0000;
	mem[2196] = 4'b0000;
	mem[2197] = 4'b0000;
	mem[2198] = 4'b0000;
	mem[2199] = 4'b0000;
	mem[2200] = 4'b0000;
	mem[2201] = 4'b0000;
	mem[2202] = 4'b0000;
	mem[2203] = 4'b0001;
	mem[2204] = 4'b0000;
	mem[2205] = 4'b0000;
	mem[2206] = 4'b0000;
	mem[2207] = 4'b0000;
	mem[2208] = 4'b0000;
	mem[2209] = 4'b0000;
	mem[2210] = 4'b0000;
	mem[2211] = 4'b0000;
	mem[2212] = 4'b0000;
	mem[2213] = 4'b0000;
	mem[2214] = 4'b0000;
	mem[2215] = 4'b0000;
	mem[2216] = 4'b0000;
	mem[2217] = 4'b0000;
	mem[2218] = 4'b0000;
	mem[2219] = 4'b0000;
	mem[2220] = 4'b0000;
	mem[2221] = 4'b0000;
	mem[2222] = 4'b0000;
	mem[2223] = 4'b0000;
	mem[2224] = 4'b0000;
	mem[2225] = 4'b0000;
	mem[2226] = 4'b0000;
	mem[2227] = 4'b0000;
	mem[2228] = 4'b0000;
	mem[2229] = 4'b0000;
	mem[2230] = 4'b0000;
	mem[2231] = 4'b0000;
	mem[2232] = 4'b0000;
	mem[2233] = 4'b0000;
	mem[2234] = 4'b0000;
	mem[2235] = 4'b0000;
	mem[2236] = 4'b0000;
	mem[2237] = 4'b0000;
	mem[2238] = 4'b0001;
	mem[2239] = 4'b0000;
	mem[2240] = 4'b0000;
	mem[2241] = 4'b0000;
	mem[2242] = 4'b0000;
	mem[2243] = 4'b0000;
	mem[2244] = 4'b0000;
	mem[2245] = 4'b0000;
	mem[2246] = 4'b0000;
	mem[2247] = 4'b0000;
	mem[2248] = 4'b0000;
	mem[2249] = 4'b0000;
	mem[2250] = 4'b0000;
	mem[2251] = 4'b0000;
	mem[2252] = 4'b0000;
	mem[2253] = 4'b0000;
	mem[2254] = 4'b0000;
	mem[2255] = 4'b0000;
	mem[2256] = 4'b0000;
	mem[2257] = 4'b0000;
	mem[2258] = 4'b0000;
	mem[2259] = 4'b0000;
	mem[2260] = 4'b0000;
	mem[2261] = 4'b0000;
	mem[2262] = 4'b0000;
	mem[2263] = 4'b0000;
	mem[2264] = 4'b0000;
	mem[2265] = 4'b0000;
	mem[2266] = 4'b0000;
	mem[2267] = 4'b0000;
	mem[2268] = 4'b0000;
	mem[2269] = 4'b0000;
	mem[2270] = 4'b0000;
	mem[2271] = 4'b0000;
	mem[2272] = 4'b0000;
	mem[2273] = 4'b0000;
	mem[2274] = 4'b0000;
	mem[2275] = 4'b0000;
	mem[2276] = 4'b0000;
	mem[2277] = 4'b0000;
	mem[2278] = 4'b0000;
	mem[2279] = 4'b0000;
	mem[2280] = 4'b0000;
	mem[2281] = 4'b0000;
	mem[2282] = 4'b0000;
	mem[2283] = 4'b0000;
	mem[2284] = 4'b0000;
	mem[2285] = 4'b0000;
	mem[2286] = 4'b0000;
	mem[2287] = 4'b0000;
	mem[2288] = 4'b0000;
	mem[2289] = 4'b0000;
	mem[2290] = 4'b0000;
	mem[2291] = 4'b0000;
	mem[2292] = 4'b0000;
	mem[2293] = 4'b0000;
	mem[2294] = 4'b0000;
	mem[2295] = 4'b0000;
	mem[2296] = 4'b0000;
	mem[2297] = 4'b0000;
	mem[2298] = 4'b0000;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0000;
	mem[2308] = 4'b0000;
	mem[2309] = 4'b0000;
	mem[2310] = 4'b0000;
	mem[2311] = 4'b0000;
	mem[2312] = 4'b0000;
	mem[2313] = 4'b0000;
	mem[2314] = 4'b0000;
	mem[2315] = 4'b0000;
	mem[2316] = 4'b0000;
	mem[2317] = 4'b0000;
	mem[2318] = 4'b0000;
	mem[2319] = 4'b0000;
	mem[2320] = 4'b0000;
	mem[2321] = 4'b0000;
	mem[2322] = 4'b0000;
	mem[2323] = 4'b0000;
	mem[2324] = 4'b0000;
	mem[2325] = 4'b0000;
	mem[2326] = 4'b0000;
	mem[2327] = 4'b0000;
	mem[2328] = 4'b0000;
	mem[2329] = 4'b0000;
	mem[2330] = 4'b0001;
	mem[2331] = 4'b0001;
	mem[2332] = 4'b0000;
	mem[2333] = 4'b0000;
	mem[2334] = 4'b0000;
	mem[2335] = 4'b0000;
	mem[2336] = 4'b0000;
	mem[2337] = 4'b0000;
	mem[2338] = 4'b0000;
	mem[2339] = 4'b0000;
	mem[2340] = 4'b0000;
	mem[2341] = 4'b0000;
	mem[2342] = 4'b0000;
	mem[2343] = 4'b0000;
	mem[2344] = 4'b0000;
	mem[2345] = 4'b0000;
	mem[2346] = 4'b0000;
	mem[2347] = 4'b0000;
	mem[2348] = 4'b0000;
	mem[2349] = 4'b0000;
	mem[2350] = 4'b0000;
	mem[2351] = 4'b0000;
	mem[2352] = 4'b0000;
	mem[2353] = 4'b0000;
	mem[2354] = 4'b0000;
	mem[2355] = 4'b0000;
	mem[2356] = 4'b0000;
	mem[2357] = 4'b0000;
	mem[2358] = 4'b0000;
	mem[2359] = 4'b0000;
	mem[2360] = 4'b0000;
	mem[2361] = 4'b0000;
	mem[2362] = 4'b0000;
	mem[2363] = 4'b0000;
	mem[2364] = 4'b0000;
	mem[2365] = 4'b0000;
	mem[2366] = 4'b0000;
	mem[2367] = 4'b0000;
	mem[2368] = 4'b0000;
	mem[2369] = 4'b0000;
	mem[2370] = 4'b0000;
	mem[2371] = 4'b0000;
	mem[2372] = 4'b0001;
	mem[2373] = 4'b0000;
	mem[2374] = 4'b0000;
	mem[2375] = 4'b0000;
	mem[2376] = 4'b0000;
	mem[2377] = 4'b0000;
	mem[2378] = 4'b0000;
	mem[2379] = 4'b0000;
	mem[2380] = 4'b0000;
	mem[2381] = 4'b0000;
	mem[2382] = 4'b0000;
	mem[2383] = 4'b0000;
	mem[2384] = 4'b0000;
	mem[2385] = 4'b0000;
	mem[2386] = 4'b0000;
	mem[2387] = 4'b0000;
	mem[2388] = 4'b0000;
	mem[2389] = 4'b0000;
	mem[2390] = 4'b0000;
	mem[2391] = 4'b0000;
	mem[2392] = 4'b0000;
	mem[2393] = 4'b0000;
	mem[2394] = 4'b0000;
	mem[2395] = 4'b0000;
	mem[2396] = 4'b0000;
	mem[2397] = 4'b0000;
	mem[2398] = 4'b0000;
	mem[2399] = 4'b0000;
	mem[2400] = 4'b0000;
	mem[2401] = 4'b0000;
	mem[2402] = 4'b0000;
	mem[2403] = 4'b0000;
	mem[2404] = 4'b0000;
	mem[2405] = 4'b0000;
	mem[2406] = 4'b0000;
	mem[2407] = 4'b0000;
	mem[2408] = 4'b0000;
	mem[2409] = 4'b0000;
	mem[2410] = 4'b0000;
	mem[2411] = 4'b0000;
	mem[2412] = 4'b0000;
	mem[2413] = 4'b0000;
	mem[2414] = 4'b0000;
	mem[2415] = 4'b0000;
	mem[2416] = 4'b0000;
	mem[2417] = 4'b0000;
	mem[2418] = 4'b0000;
	mem[2419] = 4'b0000;
	mem[2420] = 4'b0000;
	mem[2421] = 4'b0000;
	mem[2422] = 4'b0000;
	mem[2423] = 4'b0000;
	mem[2424] = 4'b0000;
	mem[2425] = 4'b0000;
	mem[2426] = 4'b0000;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0000;
	mem[2436] = 4'b0000;
	mem[2437] = 4'b0000;
	mem[2438] = 4'b0000;
	mem[2439] = 4'b0000;
	mem[2440] = 4'b0000;
	mem[2441] = 4'b0000;
	mem[2442] = 4'b0000;
	mem[2443] = 4'b0000;
	mem[2444] = 4'b0000;
	mem[2445] = 4'b0000;
	mem[2446] = 4'b0000;
	mem[2447] = 4'b0000;
	mem[2448] = 4'b0000;
	mem[2449] = 4'b0000;
	mem[2450] = 4'b0000;
	mem[2451] = 4'b0000;
	mem[2452] = 4'b0000;
	mem[2453] = 4'b0000;
	mem[2454] = 4'b0000;
	mem[2455] = 4'b0000;
	mem[2456] = 4'b0000;
	mem[2457] = 4'b0001;
	mem[2458] = 4'b0001;
	mem[2459] = 4'b0000;
	mem[2460] = 4'b0000;
	mem[2461] = 4'b0000;
	mem[2462] = 4'b0000;
	mem[2463] = 4'b0000;
	mem[2464] = 4'b0000;
	mem[2465] = 4'b0000;
	mem[2466] = 4'b0000;
	mem[2467] = 4'b0000;
	mem[2468] = 4'b0000;
	mem[2469] = 4'b0000;
	mem[2470] = 4'b0000;
	mem[2471] = 4'b0000;
	mem[2472] = 4'b0000;
	mem[2473] = 4'b0000;
	mem[2474] = 4'b0000;
	mem[2475] = 4'b0000;
	mem[2476] = 4'b0000;
	mem[2477] = 4'b0000;
	mem[2478] = 4'b0000;
	mem[2479] = 4'b0000;
	mem[2480] = 4'b0000;
	mem[2481] = 4'b0000;
	mem[2482] = 4'b0000;
	mem[2483] = 4'b0000;
	mem[2484] = 4'b0000;
	mem[2485] = 4'b0000;
	mem[2486] = 4'b0000;
	mem[2487] = 4'b0000;
	mem[2488] = 4'b0000;
	mem[2489] = 4'b0000;
	mem[2490] = 4'b0000;
	mem[2491] = 4'b0000;
	mem[2492] = 4'b0000;
	mem[2493] = 4'b0000;
	mem[2494] = 4'b0000;
	mem[2495] = 4'b0000;
	mem[2496] = 4'b0000;
	mem[2497] = 4'b0000;
	mem[2498] = 4'b0000;
	mem[2499] = 4'b0000;
	mem[2500] = 4'b0001;
	mem[2501] = 4'b0000;
	mem[2502] = 4'b0000;
	mem[2503] = 4'b0000;
	mem[2504] = 4'b0000;
	mem[2505] = 4'b0000;
	mem[2506] = 4'b0000;
	mem[2507] = 4'b0000;
	mem[2508] = 4'b0000;
	mem[2509] = 4'b0000;
	mem[2510] = 4'b0000;
	mem[2511] = 4'b0000;
	mem[2512] = 4'b0000;
	mem[2513] = 4'b0000;
	mem[2514] = 4'b0000;
	mem[2515] = 4'b0000;
	mem[2516] = 4'b0000;
	mem[2517] = 4'b0000;
	mem[2518] = 4'b0000;
	mem[2519] = 4'b0000;
	mem[2520] = 4'b0000;
	mem[2521] = 4'b0000;
	mem[2522] = 4'b0000;
	mem[2523] = 4'b0000;
	mem[2524] = 4'b0000;
	mem[2525] = 4'b0000;
	mem[2526] = 4'b0000;
	mem[2527] = 4'b0000;
	mem[2528] = 4'b0000;
	mem[2529] = 4'b0000;
	mem[2530] = 4'b0000;
	mem[2531] = 4'b0000;
	mem[2532] = 4'b0000;
	mem[2533] = 4'b0000;
	mem[2534] = 4'b0000;
	mem[2535] = 4'b0000;
	mem[2536] = 4'b0000;
	mem[2537] = 4'b0000;
	mem[2538] = 4'b0000;
	mem[2539] = 4'b0000;
	mem[2540] = 4'b0000;
	mem[2541] = 4'b0000;
	mem[2542] = 4'b0000;
	mem[2543] = 4'b0000;
	mem[2544] = 4'b0000;
	mem[2545] = 4'b0000;
	mem[2546] = 4'b0000;
	mem[2547] = 4'b0000;
	mem[2548] = 4'b0000;
	mem[2549] = 4'b0000;
	mem[2550] = 4'b0000;
	mem[2551] = 4'b0000;
	mem[2552] = 4'b0000;
	mem[2553] = 4'b0000;
	mem[2554] = 4'b0000;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b0000;
	mem[2564] = 4'b0000;
	mem[2565] = 4'b0000;
	mem[2566] = 4'b0000;
	mem[2567] = 4'b0000;
	mem[2568] = 4'b0000;
	mem[2569] = 4'b0000;
	mem[2570] = 4'b0000;
	mem[2571] = 4'b0000;
	mem[2572] = 4'b0000;
	mem[2573] = 4'b0000;
	mem[2574] = 4'b0000;
	mem[2575] = 4'b0000;
	mem[2576] = 4'b0000;
	mem[2577] = 4'b0000;
	mem[2578] = 4'b0000;
	mem[2579] = 4'b0001;
	mem[2580] = 4'b0001;
	mem[2581] = 4'b0001;
	mem[2582] = 4'b0001;
	mem[2583] = 4'b0001;
	mem[2584] = 4'b0001;
	mem[2585] = 4'b0000;
	mem[2586] = 4'b0000;
	mem[2587] = 4'b0000;
	mem[2588] = 4'b0000;
	mem[2589] = 4'b0000;
	mem[2590] = 4'b0000;
	mem[2591] = 4'b0000;
	mem[2592] = 4'b0000;
	mem[2593] = 4'b0000;
	mem[2594] = 4'b0000;
	mem[2595] = 4'b0000;
	mem[2596] = 4'b0000;
	mem[2597] = 4'b0000;
	mem[2598] = 4'b0000;
	mem[2599] = 4'b0000;
	mem[2600] = 4'b0000;
	mem[2601] = 4'b0000;
	mem[2602] = 4'b0000;
	mem[2603] = 4'b0000;
	mem[2604] = 4'b0000;
	mem[2605] = 4'b0000;
	mem[2606] = 4'b0000;
	mem[2607] = 4'b0000;
	mem[2608] = 4'b0000;
	mem[2609] = 4'b0000;
	mem[2610] = 4'b0000;
	mem[2611] = 4'b0000;
	mem[2612] = 4'b0000;
	mem[2613] = 4'b0000;
	mem[2614] = 4'b0000;
	mem[2615] = 4'b0000;
	mem[2616] = 4'b0000;
	mem[2617] = 4'b0000;
	mem[2618] = 4'b0000;
	mem[2619] = 4'b0000;
	mem[2620] = 4'b0000;
	mem[2621] = 4'b0000;
	mem[2622] = 4'b0000;
	mem[2623] = 4'b0000;
	mem[2624] = 4'b0000;
	mem[2625] = 4'b0000;
	mem[2626] = 4'b0000;
	mem[2627] = 4'b0001;
	mem[2628] = 4'b0001;
	mem[2629] = 4'b0000;
	mem[2630] = 4'b0000;
	mem[2631] = 4'b0000;
	mem[2632] = 4'b0000;
	mem[2633] = 4'b0000;
	mem[2634] = 4'b0000;
	mem[2635] = 4'b0000;
	mem[2636] = 4'b0000;
	mem[2637] = 4'b0000;
	mem[2638] = 4'b0000;
	mem[2639] = 4'b0000;
	mem[2640] = 4'b0000;
	mem[2641] = 4'b0000;
	mem[2642] = 4'b0000;
	mem[2643] = 4'b0000;
	mem[2644] = 4'b0000;
	mem[2645] = 4'b0000;
	mem[2646] = 4'b0000;
	mem[2647] = 4'b0000;
	mem[2648] = 4'b0000;
	mem[2649] = 4'b0000;
	mem[2650] = 4'b0000;
	mem[2651] = 4'b0000;
	mem[2652] = 4'b0000;
	mem[2653] = 4'b0000;
	mem[2654] = 4'b0000;
	mem[2655] = 4'b0000;
	mem[2656] = 4'b0000;
	mem[2657] = 4'b0000;
	mem[2658] = 4'b0000;
	mem[2659] = 4'b0000;
	mem[2660] = 4'b0000;
	mem[2661] = 4'b0000;
	mem[2662] = 4'b0000;
	mem[2663] = 4'b0000;
	mem[2664] = 4'b0000;
	mem[2665] = 4'b0000;
	mem[2666] = 4'b0000;
	mem[2667] = 4'b0000;
	mem[2668] = 4'b0000;
	mem[2669] = 4'b0000;
	mem[2670] = 4'b0000;
	mem[2671] = 4'b0000;
	mem[2672] = 4'b0000;
	mem[2673] = 4'b0000;
	mem[2674] = 4'b0000;
	mem[2675] = 4'b0000;
	mem[2676] = 4'b0000;
	mem[2677] = 4'b0000;
	mem[2678] = 4'b0000;
	mem[2679] = 4'b0000;
	mem[2680] = 4'b0000;
	mem[2681] = 4'b0000;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b0000;
	mem[2692] = 4'b0000;
	mem[2693] = 4'b0000;
	mem[2694] = 4'b0000;
	mem[2695] = 4'b0000;
	mem[2696] = 4'b0000;
	mem[2697] = 4'b0000;
	mem[2698] = 4'b0000;
	mem[2699] = 4'b0000;
	mem[2700] = 4'b0000;
	mem[2701] = 4'b0000;
	mem[2702] = 4'b0000;
	mem[2703] = 4'b0000;
	mem[2704] = 4'b0000;
	mem[2705] = 4'b0000;
	mem[2706] = 4'b0000;
	mem[2707] = 4'b0000;
	mem[2708] = 4'b0000;
	mem[2709] = 4'b0000;
	mem[2710] = 4'b0000;
	mem[2711] = 4'b0000;
	mem[2712] = 4'b0000;
	mem[2713] = 4'b0000;
	mem[2714] = 4'b0000;
	mem[2715] = 4'b0000;
	mem[2716] = 4'b0000;
	mem[2717] = 4'b0000;
	mem[2718] = 4'b0000;
	mem[2719] = 4'b0000;
	mem[2720] = 4'b0000;
	mem[2721] = 4'b0000;
	mem[2722] = 4'b0000;
	mem[2723] = 4'b0000;
	mem[2724] = 4'b0000;
	mem[2725] = 4'b0000;
	mem[2726] = 4'b0000;
	mem[2727] = 4'b0000;
	mem[2728] = 4'b0000;
	mem[2729] = 4'b0000;
	mem[2730] = 4'b0000;
	mem[2731] = 4'b0000;
	mem[2732] = 4'b0000;
	mem[2733] = 4'b0000;
	mem[2734] = 4'b0000;
	mem[2735] = 4'b0000;
	mem[2736] = 4'b0000;
	mem[2737] = 4'b0000;
	mem[2738] = 4'b0000;
	mem[2739] = 4'b0000;
	mem[2740] = 4'b0000;
	mem[2741] = 4'b0000;
	mem[2742] = 4'b0000;
	mem[2743] = 4'b0000;
	mem[2744] = 4'b0000;
	mem[2745] = 4'b0000;
	mem[2746] = 4'b0000;
	mem[2747] = 4'b0000;
	mem[2748] = 4'b0000;
	mem[2749] = 4'b0000;
	mem[2750] = 4'b0001;
	mem[2751] = 4'b0000;
	mem[2752] = 4'b0000;
	mem[2753] = 4'b0000;
	mem[2754] = 4'b0001;
	mem[2755] = 4'b0001;
	mem[2756] = 4'b0000;
	mem[2757] = 4'b0000;
	mem[2758] = 4'b0000;
	mem[2759] = 4'b0000;
	mem[2760] = 4'b0000;
	mem[2761] = 4'b0000;
	mem[2762] = 4'b0000;
	mem[2763] = 4'b0000;
	mem[2764] = 4'b0000;
	mem[2765] = 4'b0000;
	mem[2766] = 4'b0000;
	mem[2767] = 4'b0000;
	mem[2768] = 4'b0000;
	mem[2769] = 4'b0000;
	mem[2770] = 4'b0000;
	mem[2771] = 4'b0000;
	mem[2772] = 4'b0000;
	mem[2773] = 4'b0000;
	mem[2774] = 4'b0000;
	mem[2775] = 4'b0000;
	mem[2776] = 4'b0000;
	mem[2777] = 4'b0000;
	mem[2778] = 4'b0000;
	mem[2779] = 4'b0000;
	mem[2780] = 4'b0000;
	mem[2781] = 4'b0000;
	mem[2782] = 4'b0000;
	mem[2783] = 4'b0000;
	mem[2784] = 4'b0000;
	mem[2785] = 4'b0000;
	mem[2786] = 4'b0000;
	mem[2787] = 4'b0000;
	mem[2788] = 4'b0000;
	mem[2789] = 4'b0000;
	mem[2790] = 4'b0000;
	mem[2791] = 4'b0000;
	mem[2792] = 4'b0000;
	mem[2793] = 4'b0000;
	mem[2794] = 4'b0000;
	mem[2795] = 4'b0000;
	mem[2796] = 4'b0000;
	mem[2797] = 4'b0000;
	mem[2798] = 4'b0000;
	mem[2799] = 4'b0000;
	mem[2800] = 4'b0000;
	mem[2801] = 4'b0000;
	mem[2802] = 4'b0000;
	mem[2803] = 4'b0000;
	mem[2804] = 4'b0000;
	mem[2805] = 4'b0000;
	mem[2806] = 4'b0000;
	mem[2807] = 4'b0000;
	mem[2808] = 4'b0000;
	mem[2809] = 4'b0000;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b0000;
	mem[2820] = 4'b0000;
	mem[2821] = 4'b0000;
	mem[2822] = 4'b0000;
	mem[2823] = 4'b0000;
	mem[2824] = 4'b0000;
	mem[2825] = 4'b0000;
	mem[2826] = 4'b0000;
	mem[2827] = 4'b0000;
	mem[2828] = 4'b0000;
	mem[2829] = 4'b0000;
	mem[2830] = 4'b0000;
	mem[2831] = 4'b0000;
	mem[2832] = 4'b0000;
	mem[2833] = 4'b0000;
	mem[2834] = 4'b0000;
	mem[2835] = 4'b0000;
	mem[2836] = 4'b0000;
	mem[2837] = 4'b0000;
	mem[2838] = 4'b0000;
	mem[2839] = 4'b0000;
	mem[2840] = 4'b0000;
	mem[2841] = 4'b0000;
	mem[2842] = 4'b0000;
	mem[2843] = 4'b0000;
	mem[2844] = 4'b0000;
	mem[2845] = 4'b0000;
	mem[2846] = 4'b0000;
	mem[2847] = 4'b0000;
	mem[2848] = 4'b0000;
	mem[2849] = 4'b0000;
	mem[2850] = 4'b0000;
	mem[2851] = 4'b0000;
	mem[2852] = 4'b0000;
	mem[2853] = 4'b0000;
	mem[2854] = 4'b0000;
	mem[2855] = 4'b0000;
	mem[2856] = 4'b0000;
	mem[2857] = 4'b0000;
	mem[2858] = 4'b0000;
	mem[2859] = 4'b0000;
	mem[2860] = 4'b0000;
	mem[2861] = 4'b0000;
	mem[2862] = 4'b0000;
	mem[2863] = 4'b0000;
	mem[2864] = 4'b0000;
	mem[2865] = 4'b0000;
	mem[2866] = 4'b0000;
	mem[2867] = 4'b0000;
	mem[2868] = 4'b0000;
	mem[2869] = 4'b0000;
	mem[2870] = 4'b0000;
	mem[2871] = 4'b0000;
	mem[2872] = 4'b0000;
	mem[2873] = 4'b0000;
	mem[2874] = 4'b0000;
	mem[2875] = 4'b0000;
	mem[2876] = 4'b0000;
	mem[2877] = 4'b0000;
	mem[2878] = 4'b0000;
	mem[2879] = 4'b0000;
	mem[2880] = 4'b0001;
	mem[2881] = 4'b0001;
	mem[2882] = 4'b0000;
	mem[2883] = 4'b0000;
	mem[2884] = 4'b0000;
	mem[2885] = 4'b0000;
	mem[2886] = 4'b0000;
	mem[2887] = 4'b0000;
	mem[2888] = 4'b0000;
	mem[2889] = 4'b0000;
	mem[2890] = 4'b0000;
	mem[2891] = 4'b0000;
	mem[2892] = 4'b0000;
	mem[2893] = 4'b0000;
	mem[2894] = 4'b0000;
	mem[2895] = 4'b0000;
	mem[2896] = 4'b0000;
	mem[2897] = 4'b0000;
	mem[2898] = 4'b0000;
	mem[2899] = 4'b0000;
	mem[2900] = 4'b0000;
	mem[2901] = 4'b0000;
	mem[2902] = 4'b0000;
	mem[2903] = 4'b0000;
	mem[2904] = 4'b0000;
	mem[2905] = 4'b0000;
	mem[2906] = 4'b0000;
	mem[2907] = 4'b0000;
	mem[2908] = 4'b0000;
	mem[2909] = 4'b0000;
	mem[2910] = 4'b0000;
	mem[2911] = 4'b0000;
	mem[2912] = 4'b0000;
	mem[2913] = 4'b0000;
	mem[2914] = 4'b0000;
	mem[2915] = 4'b0000;
	mem[2916] = 4'b0000;
	mem[2917] = 4'b0000;
	mem[2918] = 4'b0000;
	mem[2919] = 4'b0000;
	mem[2920] = 4'b0000;
	mem[2921] = 4'b0000;
	mem[2922] = 4'b0000;
	mem[2923] = 4'b0000;
	mem[2924] = 4'b0000;
	mem[2925] = 4'b0000;
	mem[2926] = 4'b0000;
	mem[2927] = 4'b0000;
	mem[2928] = 4'b0000;
	mem[2929] = 4'b0000;
	mem[2930] = 4'b0000;
	mem[2931] = 4'b0000;
	mem[2932] = 4'b0000;
	mem[2933] = 4'b0000;
	mem[2934] = 4'b0000;
	mem[2935] = 4'b0000;
	mem[2936] = 4'b0000;
	mem[2937] = 4'b0000;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b0000;
	mem[2948] = 4'b0000;
	mem[2949] = 4'b0000;
	mem[2950] = 4'b0000;
	mem[2951] = 4'b0000;
	mem[2952] = 4'b0000;
	mem[2953] = 4'b0000;
	mem[2954] = 4'b0000;
	mem[2955] = 4'b0000;
	mem[2956] = 4'b0000;
	mem[2957] = 4'b0000;
	mem[2958] = 4'b0000;
	mem[2959] = 4'b0000;
	mem[2960] = 4'b0000;
	mem[2961] = 4'b0000;
	mem[2962] = 4'b0000;
	mem[2963] = 4'b0000;
	mem[2964] = 4'b0000;
	mem[2965] = 4'b0000;
	mem[2966] = 4'b0000;
	mem[2967] = 4'b0000;
	mem[2968] = 4'b0000;
	mem[2969] = 4'b0000;
	mem[2970] = 4'b0000;
	mem[2971] = 4'b0000;
	mem[2972] = 4'b0000;
	mem[2973] = 4'b0000;
	mem[2974] = 4'b0000;
	mem[2975] = 4'b0000;
	mem[2976] = 4'b0000;
	mem[2977] = 4'b0000;
	mem[2978] = 4'b0000;
	mem[2979] = 4'b0000;
	mem[2980] = 4'b0000;
	mem[2981] = 4'b0000;
	mem[2982] = 4'b0000;
	mem[2983] = 4'b0000;
	mem[2984] = 4'b0000;
	mem[2985] = 4'b0000;
	mem[2986] = 4'b0000;
	mem[2987] = 4'b0000;
	mem[2988] = 4'b0000;
	mem[2989] = 4'b0000;
	mem[2990] = 4'b0000;
	mem[2991] = 4'b0000;
	mem[2992] = 4'b0000;
	mem[2993] = 4'b0000;
	mem[2994] = 4'b0000;
	mem[2995] = 4'b0000;
	mem[2996] = 4'b0000;
	mem[2997] = 4'b0000;
	mem[2998] = 4'b0000;
	mem[2999] = 4'b0000;
	mem[3000] = 4'b0000;
	mem[3001] = 4'b0000;
	mem[3002] = 4'b0000;
	mem[3003] = 4'b0000;
	mem[3004] = 4'b0000;
	mem[3005] = 4'b0000;
	mem[3006] = 4'b0000;
	mem[3007] = 4'b0000;
	mem[3008] = 4'b0000;
	mem[3009] = 4'b0000;
	mem[3010] = 4'b0000;
	mem[3011] = 4'b0000;
	mem[3012] = 4'b0000;
	mem[3013] = 4'b0000;
	mem[3014] = 4'b0000;
	mem[3015] = 4'b0000;
	mem[3016] = 4'b0000;
	mem[3017] = 4'b0000;
	mem[3018] = 4'b0000;
	mem[3019] = 4'b0000;
	mem[3020] = 4'b0000;
	mem[3021] = 4'b0000;
	mem[3022] = 4'b0000;
	mem[3023] = 4'b0000;
	mem[3024] = 4'b0000;
	mem[3025] = 4'b0000;
	mem[3026] = 4'b0000;
	mem[3027] = 4'b0000;
	mem[3028] = 4'b0000;
	mem[3029] = 4'b0000;
	mem[3030] = 4'b0000;
	mem[3031] = 4'b0000;
	mem[3032] = 4'b0000;
	mem[3033] = 4'b0000;
	mem[3034] = 4'b0000;
	mem[3035] = 4'b0000;
	mem[3036] = 4'b0000;
	mem[3037] = 4'b0000;
	mem[3038] = 4'b0000;
	mem[3039] = 4'b0000;
	mem[3040] = 4'b0000;
	mem[3041] = 4'b0000;
	mem[3042] = 4'b0000;
	mem[3043] = 4'b0000;
	mem[3044] = 4'b0000;
	mem[3045] = 4'b0000;
	mem[3046] = 4'b0000;
	mem[3047] = 4'b0000;
	mem[3048] = 4'b0000;
	mem[3049] = 4'b0000;
	mem[3050] = 4'b0000;
	mem[3051] = 4'b0000;
	mem[3052] = 4'b0000;
	mem[3053] = 4'b0000;
	mem[3054] = 4'b0000;
	mem[3055] = 4'b0000;
	mem[3056] = 4'b0000;
	mem[3057] = 4'b0000;
	mem[3058] = 4'b0000;
	mem[3059] = 4'b0000;
	mem[3060] = 4'b0000;
	mem[3061] = 4'b0000;
	mem[3062] = 4'b0000;
	mem[3063] = 4'b0000;
	mem[3064] = 4'b0000;
	mem[3065] = 4'b0000;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b0000;
	mem[3076] = 4'b0000;
	mem[3077] = 4'b0000;
	mem[3078] = 4'b0000;
	mem[3079] = 4'b0000;
	mem[3080] = 4'b0000;
	mem[3081] = 4'b0000;
	mem[3082] = 4'b0000;
	mem[3083] = 4'b0000;
	mem[3084] = 4'b0000;
	mem[3085] = 4'b0000;
	mem[3086] = 4'b0000;
	mem[3087] = 4'b0000;
	mem[3088] = 4'b0000;
	mem[3089] = 4'b0000;
	mem[3090] = 4'b0000;
	mem[3091] = 4'b0000;
	mem[3092] = 4'b0000;
	mem[3093] = 4'b0000;
	mem[3094] = 4'b0000;
	mem[3095] = 4'b0000;
	mem[3096] = 4'b0000;
	mem[3097] = 4'b0000;
	mem[3098] = 4'b0000;
	mem[3099] = 4'b0000;
	mem[3100] = 4'b0000;
	mem[3101] = 4'b0000;
	mem[3102] = 4'b0000;
	mem[3103] = 4'b0000;
	mem[3104] = 4'b0000;
	mem[3105] = 4'b0000;
	mem[3106] = 4'b0000;
	mem[3107] = 4'b0000;
	mem[3108] = 4'b0000;
	mem[3109] = 4'b0000;
	mem[3110] = 4'b0000;
	mem[3111] = 4'b0000;
	mem[3112] = 4'b0000;
	mem[3113] = 4'b0000;
	mem[3114] = 4'b0000;
	mem[3115] = 4'b0000;
	mem[3116] = 4'b0000;
	mem[3117] = 4'b0000;
	mem[3118] = 4'b0000;
	mem[3119] = 4'b0000;
	mem[3120] = 4'b0000;
	mem[3121] = 4'b0000;
	mem[3122] = 4'b0000;
	mem[3123] = 4'b0000;
	mem[3124] = 4'b0000;
	mem[3125] = 4'b0000;
	mem[3126] = 4'b0000;
	mem[3127] = 4'b0000;
	mem[3128] = 4'b0000;
	mem[3129] = 4'b0000;
	mem[3130] = 4'b0000;
	mem[3131] = 4'b0000;
	mem[3132] = 4'b0000;
	mem[3133] = 4'b0000;
	mem[3134] = 4'b0000;
	mem[3135] = 4'b0000;
	mem[3136] = 4'b0000;
	mem[3137] = 4'b0000;
	mem[3138] = 4'b0000;
	mem[3139] = 4'b0000;
	mem[3140] = 4'b0000;
	mem[3141] = 4'b0000;
	mem[3142] = 4'b0000;
	mem[3143] = 4'b0000;
	mem[3144] = 4'b0000;
	mem[3145] = 4'b0000;
	mem[3146] = 4'b0000;
	mem[3147] = 4'b0000;
	mem[3148] = 4'b0000;
	mem[3149] = 4'b0000;
	mem[3150] = 4'b0000;
	mem[3151] = 4'b0000;
	mem[3152] = 4'b0000;
	mem[3153] = 4'b0000;
	mem[3154] = 4'b0000;
	mem[3155] = 4'b0000;
	mem[3156] = 4'b0000;
	mem[3157] = 4'b0000;
	mem[3158] = 4'b0000;
	mem[3159] = 4'b0000;
	mem[3160] = 4'b0000;
	mem[3161] = 4'b0000;
	mem[3162] = 4'b0000;
	mem[3163] = 4'b0000;
	mem[3164] = 4'b0000;
	mem[3165] = 4'b0000;
	mem[3166] = 4'b0000;
	mem[3167] = 4'b0000;
	mem[3168] = 4'b0000;
	mem[3169] = 4'b0000;
	mem[3170] = 4'b0000;
	mem[3171] = 4'b0000;
	mem[3172] = 4'b0000;
	mem[3173] = 4'b0000;
	mem[3174] = 4'b0000;
	mem[3175] = 4'b0000;
	mem[3176] = 4'b0000;
	mem[3177] = 4'b0000;
	mem[3178] = 4'b0000;
	mem[3179] = 4'b0000;
	mem[3180] = 4'b0000;
	mem[3181] = 4'b0000;
	mem[3182] = 4'b0000;
	mem[3183] = 4'b0000;
	mem[3184] = 4'b0000;
	mem[3185] = 4'b0000;
	mem[3186] = 4'b0000;
	mem[3187] = 4'b0000;
	mem[3188] = 4'b0000;
	mem[3189] = 4'b0000;
	mem[3190] = 4'b0000;
	mem[3191] = 4'b0000;
	mem[3192] = 4'b0000;
	mem[3193] = 4'b0000;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b0000;
	mem[3204] = 4'b0000;
	mem[3205] = 4'b0000;
	mem[3206] = 4'b0000;
	mem[3207] = 4'b0000;
	mem[3208] = 4'b0000;
	mem[3209] = 4'b0000;
	mem[3210] = 4'b0000;
	mem[3211] = 4'b0000;
	mem[3212] = 4'b0000;
	mem[3213] = 4'b0000;
	mem[3214] = 4'b0000;
	mem[3215] = 4'b0000;
	mem[3216] = 4'b0000;
	mem[3217] = 4'b0000;
	mem[3218] = 4'b0000;
	mem[3219] = 4'b0000;
	mem[3220] = 4'b0000;
	mem[3221] = 4'b0000;
	mem[3222] = 4'b0000;
	mem[3223] = 4'b0000;
	mem[3224] = 4'b0000;
	mem[3225] = 4'b0000;
	mem[3226] = 4'b0000;
	mem[3227] = 4'b0000;
	mem[3228] = 4'b0000;
	mem[3229] = 4'b0000;
	mem[3230] = 4'b0000;
	mem[3231] = 4'b0000;
	mem[3232] = 4'b0000;
	mem[3233] = 4'b0000;
	mem[3234] = 4'b0000;
	mem[3235] = 4'b0000;
	mem[3236] = 4'b0000;
	mem[3237] = 4'b0000;
	mem[3238] = 4'b0000;
	mem[3239] = 4'b0000;
	mem[3240] = 4'b0000;
	mem[3241] = 4'b0000;
	mem[3242] = 4'b0000;
	mem[3243] = 4'b0000;
	mem[3244] = 4'b0000;
	mem[3245] = 4'b0000;
	mem[3246] = 4'b0000;
	mem[3247] = 4'b0000;
	mem[3248] = 4'b0000;
	mem[3249] = 4'b0000;
	mem[3250] = 4'b0000;
	mem[3251] = 4'b0000;
	mem[3252] = 4'b0000;
	mem[3253] = 4'b0000;
	mem[3254] = 4'b0000;
	mem[3255] = 4'b0000;
	mem[3256] = 4'b0000;
	mem[3257] = 4'b0000;
	mem[3258] = 4'b0000;
	mem[3259] = 4'b0000;
	mem[3260] = 4'b0000;
	mem[3261] = 4'b0000;
	mem[3262] = 4'b0001;
	mem[3263] = 4'b0000;
	mem[3264] = 4'b0000;
	mem[3265] = 4'b0000;
	mem[3266] = 4'b0000;
	mem[3267] = 4'b0000;
	mem[3268] = 4'b0000;
	mem[3269] = 4'b0000;
	mem[3270] = 4'b0000;
	mem[3271] = 4'b0000;
	mem[3272] = 4'b0000;
	mem[3273] = 4'b0000;
	mem[3274] = 4'b0000;
	mem[3275] = 4'b0000;
	mem[3276] = 4'b0000;
	mem[3277] = 4'b0000;
	mem[3278] = 4'b0000;
	mem[3279] = 4'b0000;
	mem[3280] = 4'b0000;
	mem[3281] = 4'b0000;
	mem[3282] = 4'b0000;
	mem[3283] = 4'b0000;
	mem[3284] = 4'b0000;
	mem[3285] = 4'b0000;
	mem[3286] = 4'b0000;
	mem[3287] = 4'b0000;
	mem[3288] = 4'b0000;
	mem[3289] = 4'b0000;
	mem[3290] = 4'b0000;
	mem[3291] = 4'b0000;
	mem[3292] = 4'b0000;
	mem[3293] = 4'b0000;
	mem[3294] = 4'b0000;
	mem[3295] = 4'b0000;
	mem[3296] = 4'b0000;
	mem[3297] = 4'b0000;
	mem[3298] = 4'b0000;
	mem[3299] = 4'b0000;
	mem[3300] = 4'b0000;
	mem[3301] = 4'b0000;
	mem[3302] = 4'b0000;
	mem[3303] = 4'b0000;
	mem[3304] = 4'b0000;
	mem[3305] = 4'b0000;
	mem[3306] = 4'b0000;
	mem[3307] = 4'b0000;
	mem[3308] = 4'b0000;
	mem[3309] = 4'b0000;
	mem[3310] = 4'b0000;
	mem[3311] = 4'b0000;
	mem[3312] = 4'b0000;
	mem[3313] = 4'b0000;
	mem[3314] = 4'b0000;
	mem[3315] = 4'b0000;
	mem[3316] = 4'b0000;
	mem[3317] = 4'b0000;
	mem[3318] = 4'b0000;
	mem[3319] = 4'b0000;
	mem[3320] = 4'b0000;
	mem[3321] = 4'b0000;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b0000;
	mem[3332] = 4'b0000;
	mem[3333] = 4'b0000;
	mem[3334] = 4'b0000;
	mem[3335] = 4'b0000;
	mem[3336] = 4'b0000;
	mem[3337] = 4'b0000;
	mem[3338] = 4'b0000;
	mem[3339] = 4'b0000;
	mem[3340] = 4'b0000;
	mem[3341] = 4'b0000;
	mem[3342] = 4'b0000;
	mem[3343] = 4'b0000;
	mem[3344] = 4'b0000;
	mem[3345] = 4'b0000;
	mem[3346] = 4'b0001;
	mem[3347] = 4'b0001;
	mem[3348] = 4'b0000;
	mem[3349] = 4'b0000;
	mem[3350] = 4'b0000;
	mem[3351] = 4'b0000;
	mem[3352] = 4'b0000;
	mem[3353] = 4'b0000;
	mem[3354] = 4'b0000;
	mem[3355] = 4'b0000;
	mem[3356] = 4'b0000;
	mem[3357] = 4'b0000;
	mem[3358] = 4'b0000;
	mem[3359] = 4'b0000;
	mem[3360] = 4'b0000;
	mem[3361] = 4'b0000;
	mem[3362] = 4'b0000;
	mem[3363] = 4'b0000;
	mem[3364] = 4'b0000;
	mem[3365] = 4'b0000;
	mem[3366] = 4'b0000;
	mem[3367] = 4'b0000;
	mem[3368] = 4'b0000;
	mem[3369] = 4'b0000;
	mem[3370] = 4'b0000;
	mem[3371] = 4'b0000;
	mem[3372] = 4'b0000;
	mem[3373] = 4'b0000;
	mem[3374] = 4'b0000;
	mem[3375] = 4'b0000;
	mem[3376] = 4'b0000;
	mem[3377] = 4'b0000;
	mem[3378] = 4'b0000;
	mem[3379] = 4'b0000;
	mem[3380] = 4'b0000;
	mem[3381] = 4'b0000;
	mem[3382] = 4'b0000;
	mem[3383] = 4'b0000;
	mem[3384] = 4'b0000;
	mem[3385] = 4'b0000;
	mem[3386] = 4'b0000;
	mem[3387] = 4'b0000;
	mem[3388] = 4'b0000;
	mem[3389] = 4'b0001;
	mem[3390] = 4'b0001;
	mem[3391] = 4'b0000;
	mem[3392] = 4'b0000;
	mem[3393] = 4'b0000;
	mem[3394] = 4'b0000;
	mem[3395] = 4'b0000;
	mem[3396] = 4'b0000;
	mem[3397] = 4'b0000;
	mem[3398] = 4'b0000;
	mem[3399] = 4'b0000;
	mem[3400] = 4'b0000;
	mem[3401] = 4'b0000;
	mem[3402] = 4'b0000;
	mem[3403] = 4'b0000;
	mem[3404] = 4'b0000;
	mem[3405] = 4'b0000;
	mem[3406] = 4'b0000;
	mem[3407] = 4'b0000;
	mem[3408] = 4'b0000;
	mem[3409] = 4'b0000;
	mem[3410] = 4'b0000;
	mem[3411] = 4'b0000;
	mem[3412] = 4'b0000;
	mem[3413] = 4'b0000;
	mem[3414] = 4'b0000;
	mem[3415] = 4'b0000;
	mem[3416] = 4'b0000;
	mem[3417] = 4'b0000;
	mem[3418] = 4'b0000;
	mem[3419] = 4'b0000;
	mem[3420] = 4'b0000;
	mem[3421] = 4'b0000;
	mem[3422] = 4'b0000;
	mem[3423] = 4'b0000;
	mem[3424] = 4'b0000;
	mem[3425] = 4'b0000;
	mem[3426] = 4'b0000;
	mem[3427] = 4'b0000;
	mem[3428] = 4'b0000;
	mem[3429] = 4'b0000;
	mem[3430] = 4'b0000;
	mem[3431] = 4'b0000;
	mem[3432] = 4'b0000;
	mem[3433] = 4'b0000;
	mem[3434] = 4'b0000;
	mem[3435] = 4'b0000;
	mem[3436] = 4'b0000;
	mem[3437] = 4'b0000;
	mem[3438] = 4'b0000;
	mem[3439] = 4'b0000;
	mem[3440] = 4'b0000;
	mem[3441] = 4'b0000;
	mem[3442] = 4'b0000;
	mem[3443] = 4'b0000;
	mem[3444] = 4'b0000;
	mem[3445] = 4'b0000;
	mem[3446] = 4'b0000;
	mem[3447] = 4'b0000;
	mem[3448] = 4'b0000;
	mem[3449] = 4'b0000;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b0000;
	mem[3460] = 4'b0000;
	mem[3461] = 4'b0000;
	mem[3462] = 4'b0000;
	mem[3463] = 4'b0000;
	mem[3464] = 4'b0000;
	mem[3465] = 4'b0000;
	mem[3466] = 4'b0000;
	mem[3467] = 4'b0000;
	mem[3468] = 4'b0000;
	mem[3469] = 4'b0000;
	mem[3470] = 4'b0000;
	mem[3471] = 4'b0000;
	mem[3472] = 4'b0000;
	mem[3473] = 4'b0001;
	mem[3474] = 4'b0001;
	mem[3475] = 4'b0000;
	mem[3476] = 4'b0000;
	mem[3477] = 4'b0000;
	mem[3478] = 4'b0000;
	mem[3479] = 4'b0000;
	mem[3480] = 4'b0000;
	mem[3481] = 4'b0000;
	mem[3482] = 4'b0000;
	mem[3483] = 4'b0000;
	mem[3484] = 4'b0000;
	mem[3485] = 4'b0000;
	mem[3486] = 4'b0000;
	mem[3487] = 4'b0000;
	mem[3488] = 4'b0000;
	mem[3489] = 4'b0000;
	mem[3490] = 4'b0000;
	mem[3491] = 4'b0000;
	mem[3492] = 4'b0000;
	mem[3493] = 4'b0000;
	mem[3494] = 4'b0000;
	mem[3495] = 4'b0000;
	mem[3496] = 4'b0000;
	mem[3497] = 4'b0000;
	mem[3498] = 4'b0000;
	mem[3499] = 4'b0000;
	mem[3500] = 4'b0000;
	mem[3501] = 4'b0000;
	mem[3502] = 4'b0000;
	mem[3503] = 4'b0000;
	mem[3504] = 4'b0000;
	mem[3505] = 4'b0000;
	mem[3506] = 4'b0000;
	mem[3507] = 4'b0000;
	mem[3508] = 4'b0000;
	mem[3509] = 4'b0000;
	mem[3510] = 4'b0000;
	mem[3511] = 4'b0000;
	mem[3512] = 4'b0000;
	mem[3513] = 4'b0000;
	mem[3514] = 4'b0000;
	mem[3515] = 4'b0000;
	mem[3516] = 4'b0000;
	mem[3517] = 4'b0000;
	mem[3518] = 4'b0000;
	mem[3519] = 4'b0000;
	mem[3520] = 4'b0000;
	mem[3521] = 4'b0000;
	mem[3522] = 4'b0000;
	mem[3523] = 4'b0000;
	mem[3524] = 4'b0000;
	mem[3525] = 4'b0000;
	mem[3526] = 4'b0000;
	mem[3527] = 4'b0000;
	mem[3528] = 4'b0000;
	mem[3529] = 4'b0000;
	mem[3530] = 4'b0000;
	mem[3531] = 4'b0000;
	mem[3532] = 4'b0000;
	mem[3533] = 4'b0000;
	mem[3534] = 4'b0000;
	mem[3535] = 4'b0000;
	mem[3536] = 4'b0000;
	mem[3537] = 4'b0000;
	mem[3538] = 4'b0000;
	mem[3539] = 4'b0000;
	mem[3540] = 4'b0000;
	mem[3541] = 4'b0000;
	mem[3542] = 4'b0000;
	mem[3543] = 4'b0000;
	mem[3544] = 4'b0000;
	mem[3545] = 4'b0000;
	mem[3546] = 4'b0000;
	mem[3547] = 4'b0000;
	mem[3548] = 4'b0000;
	mem[3549] = 4'b0000;
	mem[3550] = 4'b0000;
	mem[3551] = 4'b0000;
	mem[3552] = 4'b0000;
	mem[3553] = 4'b0000;
	mem[3554] = 4'b0000;
	mem[3555] = 4'b0000;
	mem[3556] = 4'b0000;
	mem[3557] = 4'b0000;
	mem[3558] = 4'b0000;
	mem[3559] = 4'b0000;
	mem[3560] = 4'b0000;
	mem[3561] = 4'b0000;
	mem[3562] = 4'b0000;
	mem[3563] = 4'b0000;
	mem[3564] = 4'b0000;
	mem[3565] = 4'b0000;
	mem[3566] = 4'b0000;
	mem[3567] = 4'b0000;
	mem[3568] = 4'b0000;
	mem[3569] = 4'b0000;
	mem[3570] = 4'b0000;
	mem[3571] = 4'b0000;
	mem[3572] = 4'b0000;
	mem[3573] = 4'b0000;
	mem[3574] = 4'b0000;
	mem[3575] = 4'b0000;
	mem[3576] = 4'b0000;
	mem[3577] = 4'b0000;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b0000;
	mem[3588] = 4'b0000;
	mem[3589] = 4'b0000;
	mem[3590] = 4'b0000;
	mem[3591] = 4'b0000;
	mem[3592] = 4'b0000;
	mem[3593] = 4'b0000;
	mem[3594] = 4'b0000;
	mem[3595] = 4'b0000;
	mem[3596] = 4'b0000;
	mem[3597] = 4'b0000;
	mem[3598] = 4'b0000;
	mem[3599] = 4'b0000;
	mem[3600] = 4'b0001;
	mem[3601] = 4'b0001;
	mem[3602] = 4'b0000;
	mem[3603] = 4'b0000;
	mem[3604] = 4'b0000;
	mem[3605] = 4'b0000;
	mem[3606] = 4'b0000;
	mem[3607] = 4'b0000;
	mem[3608] = 4'b0000;
	mem[3609] = 4'b0000;
	mem[3610] = 4'b0000;
	mem[3611] = 4'b0000;
	mem[3612] = 4'b0000;
	mem[3613] = 4'b0000;
	mem[3614] = 4'b0000;
	mem[3615] = 4'b0000;
	mem[3616] = 4'b0000;
	mem[3617] = 4'b0000;
	mem[3618] = 4'b0000;
	mem[3619] = 4'b0000;
	mem[3620] = 4'b0000;
	mem[3621] = 4'b0000;
	mem[3622] = 4'b0000;
	mem[3623] = 4'b0000;
	mem[3624] = 4'b0000;
	mem[3625] = 4'b0000;
	mem[3626] = 4'b0000;
	mem[3627] = 4'b0000;
	mem[3628] = 4'b0000;
	mem[3629] = 4'b0000;
	mem[3630] = 4'b0000;
	mem[3631] = 4'b0000;
	mem[3632] = 4'b0000;
	mem[3633] = 4'b0000;
	mem[3634] = 4'b0000;
	mem[3635] = 4'b0000;
	mem[3636] = 4'b0000;
	mem[3637] = 4'b0000;
	mem[3638] = 4'b0000;
	mem[3639] = 4'b0000;
	mem[3640] = 4'b0000;
	mem[3641] = 4'b0000;
	mem[3642] = 4'b0000;
	mem[3643] = 4'b0000;
	mem[3644] = 4'b0000;
	mem[3645] = 4'b0000;
	mem[3646] = 4'b0000;
	mem[3647] = 4'b0000;
	mem[3648] = 4'b0000;
	mem[3649] = 4'b0000;
	mem[3650] = 4'b0000;
	mem[3651] = 4'b0000;
	mem[3652] = 4'b0000;
	mem[3653] = 4'b0000;
	mem[3654] = 4'b0000;
	mem[3655] = 4'b0000;
	mem[3656] = 4'b0000;
	mem[3657] = 4'b0000;
	mem[3658] = 4'b0000;
	mem[3659] = 4'b0000;
	mem[3660] = 4'b0000;
	mem[3661] = 4'b0000;
	mem[3662] = 4'b0000;
	mem[3663] = 4'b0000;
	mem[3664] = 4'b0000;
	mem[3665] = 4'b0000;
	mem[3666] = 4'b0000;
	mem[3667] = 4'b0000;
	mem[3668] = 4'b0000;
	mem[3669] = 4'b0000;
	mem[3670] = 4'b0000;
	mem[3671] = 4'b0000;
	mem[3672] = 4'b0000;
	mem[3673] = 4'b0000;
	mem[3674] = 4'b0000;
	mem[3675] = 4'b0000;
	mem[3676] = 4'b0000;
	mem[3677] = 4'b0000;
	mem[3678] = 4'b0000;
	mem[3679] = 4'b0000;
	mem[3680] = 4'b0000;
	mem[3681] = 4'b0000;
	mem[3682] = 4'b0000;
	mem[3683] = 4'b0000;
	mem[3684] = 4'b0000;
	mem[3685] = 4'b0000;
	mem[3686] = 4'b0000;
	mem[3687] = 4'b0000;
	mem[3688] = 4'b0000;
	mem[3689] = 4'b0000;
	mem[3690] = 4'b0000;
	mem[3691] = 4'b0000;
	mem[3692] = 4'b0000;
	mem[3693] = 4'b0000;
	mem[3694] = 4'b0000;
	mem[3695] = 4'b0000;
	mem[3696] = 4'b0000;
	mem[3697] = 4'b0000;
	mem[3698] = 4'b0000;
	mem[3699] = 4'b0000;
	mem[3700] = 4'b0000;
	mem[3701] = 4'b0000;
	mem[3702] = 4'b0000;
	mem[3703] = 4'b0000;
	mem[3704] = 4'b0000;
	mem[3705] = 4'b0000;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b0000;
	mem[3716] = 4'b0000;
	mem[3717] = 4'b0000;
	mem[3718] = 4'b0000;
	mem[3719] = 4'b0000;
	mem[3720] = 4'b0000;
	mem[3721] = 4'b0000;
	mem[3722] = 4'b0000;
	mem[3723] = 4'b0000;
	mem[3724] = 4'b0000;
	mem[3725] = 4'b0000;
	mem[3726] = 4'b0000;
	mem[3727] = 4'b0000;
	mem[3728] = 4'b0000;
	mem[3729] = 4'b0000;
	mem[3730] = 4'b0000;
	mem[3731] = 4'b0000;
	mem[3732] = 4'b0000;
	mem[3733] = 4'b0000;
	mem[3734] = 4'b0000;
	mem[3735] = 4'b0000;
	mem[3736] = 4'b0000;
	mem[3737] = 4'b0000;
	mem[3738] = 4'b0000;
	mem[3739] = 4'b0000;
	mem[3740] = 4'b0000;
	mem[3741] = 4'b0000;
	mem[3742] = 4'b0000;
	mem[3743] = 4'b0000;
	mem[3744] = 4'b0000;
	mem[3745] = 4'b0000;
	mem[3746] = 4'b0000;
	mem[3747] = 4'b0000;
	mem[3748] = 4'b0000;
	mem[3749] = 4'b0000;
	mem[3750] = 4'b0000;
	mem[3751] = 4'b0000;
	mem[3752] = 4'b0000;
	mem[3753] = 4'b0000;
	mem[3754] = 4'b0000;
	mem[3755] = 4'b0000;
	mem[3756] = 4'b0000;
	mem[3757] = 4'b0000;
	mem[3758] = 4'b0000;
	mem[3759] = 4'b0000;
	mem[3760] = 4'b0000;
	mem[3761] = 4'b0000;
	mem[3762] = 4'b0000;
	mem[3763] = 4'b0000;
	mem[3764] = 4'b0000;
	mem[3765] = 4'b0000;
	mem[3766] = 4'b0000;
	mem[3767] = 4'b0000;
	mem[3768] = 4'b0000;
	mem[3769] = 4'b0000;
	mem[3770] = 4'b0000;
	mem[3771] = 4'b0000;
	mem[3772] = 4'b0000;
	mem[3773] = 4'b0000;
	mem[3774] = 4'b0000;
	mem[3775] = 4'b0000;
	mem[3776] = 4'b0000;
	mem[3777] = 4'b0000;
	mem[3778] = 4'b0000;
	mem[3779] = 4'b0000;
	mem[3780] = 4'b0000;
	mem[3781] = 4'b0000;
	mem[3782] = 4'b0000;
	mem[3783] = 4'b0000;
	mem[3784] = 4'b0000;
	mem[3785] = 4'b0000;
	mem[3786] = 4'b0000;
	mem[3787] = 4'b0000;
	mem[3788] = 4'b0000;
	mem[3789] = 4'b0000;
	mem[3790] = 4'b0000;
	mem[3791] = 4'b0000;
	mem[3792] = 4'b0000;
	mem[3793] = 4'b0000;
	mem[3794] = 4'b0000;
	mem[3795] = 4'b0000;
	mem[3796] = 4'b0000;
	mem[3797] = 4'b0000;
	mem[3798] = 4'b0000;
	mem[3799] = 4'b0000;
	mem[3800] = 4'b0000;
	mem[3801] = 4'b0000;
	mem[3802] = 4'b0000;
	mem[3803] = 4'b0000;
	mem[3804] = 4'b0000;
	mem[3805] = 4'b0000;
	mem[3806] = 4'b0000;
	mem[3807] = 4'b0000;
	mem[3808] = 4'b0000;
	mem[3809] = 4'b0000;
	mem[3810] = 4'b0000;
	mem[3811] = 4'b0000;
	mem[3812] = 4'b0000;
	mem[3813] = 4'b0000;
	mem[3814] = 4'b0000;
	mem[3815] = 4'b0000;
	mem[3816] = 4'b0000;
	mem[3817] = 4'b0000;
	mem[3818] = 4'b0000;
	mem[3819] = 4'b0000;
	mem[3820] = 4'b0000;
	mem[3821] = 4'b0000;
	mem[3822] = 4'b0000;
	mem[3823] = 4'b0000;
	mem[3824] = 4'b0000;
	mem[3825] = 4'b0000;
	mem[3826] = 4'b0000;
	mem[3827] = 4'b0000;
	mem[3828] = 4'b0000;
	mem[3829] = 4'b0000;
	mem[3830] = 4'b0000;
	mem[3831] = 4'b0000;
	mem[3832] = 4'b0000;
	mem[3833] = 4'b0000;
	mem[3834] = 4'b0000;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b0000;
	mem[3844] = 4'b0000;
	mem[3845] = 4'b0000;
	mem[3846] = 4'b0000;
	mem[3847] = 4'b0000;
	mem[3848] = 4'b0000;
	mem[3849] = 4'b0000;
	mem[3850] = 4'b0000;
	mem[3851] = 4'b0000;
	mem[3852] = 4'b0000;
	mem[3853] = 4'b0000;
	mem[3854] = 4'b0000;
	mem[3855] = 4'b0000;
	mem[3856] = 4'b0000;
	mem[3857] = 4'b0000;
	mem[3858] = 4'b0000;
	mem[3859] = 4'b0000;
	mem[3860] = 4'b0000;
	mem[3861] = 4'b0000;
	mem[3862] = 4'b0000;
	mem[3863] = 4'b0000;
	mem[3864] = 4'b0000;
	mem[3865] = 4'b0000;
	mem[3866] = 4'b0000;
	mem[3867] = 4'b0000;
	mem[3868] = 4'b0000;
	mem[3869] = 4'b0000;
	mem[3870] = 4'b0000;
	mem[3871] = 4'b0000;
	mem[3872] = 4'b0000;
	mem[3873] = 4'b0000;
	mem[3874] = 4'b0000;
	mem[3875] = 4'b0000;
	mem[3876] = 4'b0000;
	mem[3877] = 4'b0000;
	mem[3878] = 4'b0000;
	mem[3879] = 4'b0000;
	mem[3880] = 4'b0000;
	mem[3881] = 4'b0000;
	mem[3882] = 4'b0000;
	mem[3883] = 4'b0000;
	mem[3884] = 4'b0000;
	mem[3885] = 4'b0000;
	mem[3886] = 4'b0000;
	mem[3887] = 4'b0000;
	mem[3888] = 4'b0000;
	mem[3889] = 4'b0000;
	mem[3890] = 4'b0000;
	mem[3891] = 4'b0000;
	mem[3892] = 4'b0000;
	mem[3893] = 4'b0000;
	mem[3894] = 4'b0000;
	mem[3895] = 4'b0000;
	mem[3896] = 4'b0000;
	mem[3897] = 4'b0000;
	mem[3898] = 4'b0000;
	mem[3899] = 4'b0000;
	mem[3900] = 4'b0000;
	mem[3901] = 4'b0000;
	mem[3902] = 4'b0000;
	mem[3903] = 4'b0000;
	mem[3904] = 4'b0000;
	mem[3905] = 4'b0000;
	mem[3906] = 4'b0000;
	mem[3907] = 4'b0000;
	mem[3908] = 4'b0000;
	mem[3909] = 4'b0000;
	mem[3910] = 4'b0000;
	mem[3911] = 4'b0000;
	mem[3912] = 4'b0000;
	mem[3913] = 4'b0000;
	mem[3914] = 4'b0000;
	mem[3915] = 4'b0000;
	mem[3916] = 4'b0000;
	mem[3917] = 4'b0000;
	mem[3918] = 4'b0000;
	mem[3919] = 4'b0000;
	mem[3920] = 4'b0000;
	mem[3921] = 4'b0000;
	mem[3922] = 4'b0000;
	mem[3923] = 4'b0000;
	mem[3924] = 4'b0000;
	mem[3925] = 4'b0000;
	mem[3926] = 4'b0000;
	mem[3927] = 4'b0000;
	mem[3928] = 4'b0000;
	mem[3929] = 4'b0000;
	mem[3930] = 4'b0000;
	mem[3931] = 4'b0000;
	mem[3932] = 4'b0000;
	mem[3933] = 4'b0000;
	mem[3934] = 4'b0000;
	mem[3935] = 4'b0000;
	mem[3936] = 4'b0000;
	mem[3937] = 4'b0000;
	mem[3938] = 4'b0000;
	mem[3939] = 4'b0000;
	mem[3940] = 4'b0000;
	mem[3941] = 4'b0000;
	mem[3942] = 4'b0000;
	mem[3943] = 4'b0000;
	mem[3944] = 4'b0000;
	mem[3945] = 4'b0000;
	mem[3946] = 4'b0000;
	mem[3947] = 4'b0000;
	mem[3948] = 4'b0000;
	mem[3949] = 4'b0000;
	mem[3950] = 4'b0000;
	mem[3951] = 4'b0000;
	mem[3952] = 4'b0000;
	mem[3953] = 4'b0000;
	mem[3954] = 4'b0000;
	mem[3955] = 4'b0000;
	mem[3956] = 4'b0000;
	mem[3957] = 4'b0000;
	mem[3958] = 4'b0000;
	mem[3959] = 4'b0000;
	mem[3960] = 4'b0000;
	mem[3961] = 4'b0000;
	mem[3962] = 4'b0000;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b0000;
	mem[3972] = 4'b0000;
	mem[3973] = 4'b0000;
	mem[3974] = 4'b0000;
	mem[3975] = 4'b0000;
	mem[3976] = 4'b0000;
	mem[3977] = 4'b0000;
	mem[3978] = 4'b0000;
	mem[3979] = 4'b0000;
	mem[3980] = 4'b0000;
	mem[3981] = 4'b0000;
	mem[3982] = 4'b0000;
	mem[3983] = 4'b0000;
	mem[3984] = 4'b0000;
	mem[3985] = 4'b0000;
	mem[3986] = 4'b0000;
	mem[3987] = 4'b0000;
	mem[3988] = 4'b0000;
	mem[3989] = 4'b0000;
	mem[3990] = 4'b0000;
	mem[3991] = 4'b0000;
	mem[3992] = 4'b0000;
	mem[3993] = 4'b0000;
	mem[3994] = 4'b0000;
	mem[3995] = 4'b0000;
	mem[3996] = 4'b0000;
	mem[3997] = 4'b0000;
	mem[3998] = 4'b0000;
	mem[3999] = 4'b0000;
	mem[4000] = 4'b0000;
	mem[4001] = 4'b0000;
	mem[4002] = 4'b0000;
	mem[4003] = 4'b0000;
	mem[4004] = 4'b0000;
	mem[4005] = 4'b0000;
	mem[4006] = 4'b0000;
	mem[4007] = 4'b0000;
	mem[4008] = 4'b0000;
	mem[4009] = 4'b0000;
	mem[4010] = 4'b0000;
	mem[4011] = 4'b0000;
	mem[4012] = 4'b0000;
	mem[4013] = 4'b0000;
	mem[4014] = 4'b0000;
	mem[4015] = 4'b0000;
	mem[4016] = 4'b0000;
	mem[4017] = 4'b0000;
	mem[4018] = 4'b0000;
	mem[4019] = 4'b0000;
	mem[4020] = 4'b0000;
	mem[4021] = 4'b0000;
	mem[4022] = 4'b0000;
	mem[4023] = 4'b0000;
	mem[4024] = 4'b0000;
	mem[4025] = 4'b0000;
	mem[4026] = 4'b0000;
	mem[4027] = 4'b0000;
	mem[4028] = 4'b0000;
	mem[4029] = 4'b0000;
	mem[4030] = 4'b0000;
	mem[4031] = 4'b0000;
	mem[4032] = 4'b0000;
	mem[4033] = 4'b0000;
	mem[4034] = 4'b0000;
	mem[4035] = 4'b0000;
	mem[4036] = 4'b0000;
	mem[4037] = 4'b0000;
	mem[4038] = 4'b0000;
	mem[4039] = 4'b0000;
	mem[4040] = 4'b0000;
	mem[4041] = 4'b0000;
	mem[4042] = 4'b0000;
	mem[4043] = 4'b0000;
	mem[4044] = 4'b0000;
	mem[4045] = 4'b0000;
	mem[4046] = 4'b0000;
	mem[4047] = 4'b0000;
	mem[4048] = 4'b0000;
	mem[4049] = 4'b0000;
	mem[4050] = 4'b0000;
	mem[4051] = 4'b0000;
	mem[4052] = 4'b0000;
	mem[4053] = 4'b0000;
	mem[4054] = 4'b0000;
	mem[4055] = 4'b0000;
	mem[4056] = 4'b0000;
	mem[4057] = 4'b0000;
	mem[4058] = 4'b0000;
	mem[4059] = 4'b0000;
	mem[4060] = 4'b0000;
	mem[4061] = 4'b0000;
	mem[4062] = 4'b0000;
	mem[4063] = 4'b0000;
	mem[4064] = 4'b0000;
	mem[4065] = 4'b0000;
	mem[4066] = 4'b0000;
	mem[4067] = 4'b0000;
	mem[4068] = 4'b0000;
	mem[4069] = 4'b0000;
	mem[4070] = 4'b0000;
	mem[4071] = 4'b0000;
	mem[4072] = 4'b0000;
	mem[4073] = 4'b0000;
	mem[4074] = 4'b0000;
	mem[4075] = 4'b0000;
	mem[4076] = 4'b0000;
	mem[4077] = 4'b0000;
	mem[4078] = 4'b0000;
	mem[4079] = 4'b0000;
	mem[4080] = 4'b0000;
	mem[4081] = 4'b0000;
	mem[4082] = 4'b0000;
	mem[4083] = 4'b0000;
	mem[4084] = 4'b0000;
	mem[4085] = 4'b0000;
	mem[4086] = 4'b0000;
	mem[4087] = 4'b0000;
	mem[4088] = 4'b0000;
	mem[4089] = 4'b0000;
	mem[4090] = 4'b0000;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_0g (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0000;
	mem[4] = 4'b0000;
	mem[5] = 4'b0000;
	mem[6] = 4'b0000;
	mem[7] = 4'b0000;
	mem[8] = 4'b0000;
	mem[9] = 4'b0000;
	mem[10] = 4'b0000;
	mem[11] = 4'b0000;
	mem[12] = 4'b0000;
	mem[13] = 4'b0000;
	mem[14] = 4'b0000;
	mem[15] = 4'b0000;
	mem[16] = 4'b0000;
	mem[17] = 4'b0000;
	mem[18] = 4'b0000;
	mem[19] = 4'b0000;
	mem[20] = 4'b0000;
	mem[21] = 4'b0000;
	mem[22] = 4'b0000;
	mem[23] = 4'b0000;
	mem[24] = 4'b0000;
	mem[25] = 4'b0000;
	mem[26] = 4'b0000;
	mem[27] = 4'b0000;
	mem[28] = 4'b0000;
	mem[29] = 4'b0000;
	mem[30] = 4'b0000;
	mem[31] = 4'b0000;
	mem[32] = 4'b0000;
	mem[33] = 4'b0000;
	mem[34] = 4'b0000;
	mem[35] = 4'b0000;
	mem[36] = 4'b0000;
	mem[37] = 4'b0000;
	mem[38] = 4'b0000;
	mem[39] = 4'b0000;
	mem[40] = 4'b0000;
	mem[41] = 4'b0000;
	mem[42] = 4'b0000;
	mem[43] = 4'b0000;
	mem[44] = 4'b0000;
	mem[45] = 4'b0000;
	mem[46] = 4'b0000;
	mem[47] = 4'b0000;
	mem[48] = 4'b0000;
	mem[49] = 4'b0000;
	mem[50] = 4'b0000;
	mem[51] = 4'b0000;
	mem[52] = 4'b0000;
	mem[53] = 4'b0000;
	mem[54] = 4'b0000;
	mem[55] = 4'b0000;
	mem[56] = 4'b0000;
	mem[57] = 4'b0000;
	mem[58] = 4'b0000;
	mem[59] = 4'b0000;
	mem[60] = 4'b0000;
	mem[61] = 4'b0000;
	mem[62] = 4'b0000;
	mem[63] = 4'b0000;
	mem[64] = 4'b0000;
	mem[65] = 4'b0000;
	mem[66] = 4'b0000;
	mem[67] = 4'b0000;
	mem[68] = 4'b0000;
	mem[69] = 4'b0000;
	mem[70] = 4'b0000;
	mem[71] = 4'b0000;
	mem[72] = 4'b0000;
	mem[73] = 4'b0000;
	mem[74] = 4'b0000;
	mem[75] = 4'b0000;
	mem[76] = 4'b0000;
	mem[77] = 4'b0000;
	mem[78] = 4'b0000;
	mem[79] = 4'b0000;
	mem[80] = 4'b0000;
	mem[81] = 4'b0000;
	mem[82] = 4'b0000;
	mem[83] = 4'b0000;
	mem[84] = 4'b0000;
	mem[85] = 4'b0000;
	mem[86] = 4'b0000;
	mem[87] = 4'b0000;
	mem[88] = 4'b0000;
	mem[89] = 4'b0000;
	mem[90] = 4'b0000;
	mem[91] = 4'b0000;
	mem[92] = 4'b0000;
	mem[93] = 4'b0000;
	mem[94] = 4'b0000;
	mem[95] = 4'b0000;
	mem[96] = 4'b0000;
	mem[97] = 4'b0000;
	mem[98] = 4'b0000;
	mem[99] = 4'b0000;
	mem[100] = 4'b0000;
	mem[101] = 4'b0000;
	mem[102] = 4'b0000;
	mem[103] = 4'b0000;
	mem[104] = 4'b0000;
	mem[105] = 4'b0000;
	mem[106] = 4'b0000;
	mem[107] = 4'b0000;
	mem[108] = 4'b0000;
	mem[109] = 4'b0000;
	mem[110] = 4'b0000;
	mem[111] = 4'b0000;
	mem[112] = 4'b0000;
	mem[113] = 4'b0000;
	mem[114] = 4'b0000;
	mem[115] = 4'b0000;
	mem[116] = 4'b0000;
	mem[117] = 4'b0000;
	mem[118] = 4'b0000;
	mem[119] = 4'b0000;
	mem[120] = 4'b0000;
	mem[121] = 4'b0000;
	mem[122] = 4'b0000;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b0000;
	mem[132] = 4'b0000;
	mem[133] = 4'b0000;
	mem[134] = 4'b0000;
	mem[135] = 4'b0000;
	mem[136] = 4'b0000;
	mem[137] = 4'b0000;
	mem[138] = 4'b0000;
	mem[139] = 4'b0000;
	mem[140] = 4'b0000;
	mem[141] = 4'b0000;
	mem[142] = 4'b0000;
	mem[143] = 4'b0000;
	mem[144] = 4'b0000;
	mem[145] = 4'b0000;
	mem[146] = 4'b0000;
	mem[147] = 4'b0000;
	mem[148] = 4'b0000;
	mem[149] = 4'b0000;
	mem[150] = 4'b0000;
	mem[151] = 4'b0000;
	mem[152] = 4'b0000;
	mem[153] = 4'b0000;
	mem[154] = 4'b0000;
	mem[155] = 4'b0000;
	mem[156] = 4'b0000;
	mem[157] = 4'b0000;
	mem[158] = 4'b0000;
	mem[159] = 4'b0000;
	mem[160] = 4'b0000;
	mem[161] = 4'b0000;
	mem[162] = 4'b0000;
	mem[163] = 4'b0000;
	mem[164] = 4'b0000;
	mem[165] = 4'b0000;
	mem[166] = 4'b0000;
	mem[167] = 4'b0000;
	mem[168] = 4'b0000;
	mem[169] = 4'b0000;
	mem[170] = 4'b0000;
	mem[171] = 4'b0000;
	mem[172] = 4'b0000;
	mem[173] = 4'b0000;
	mem[174] = 4'b0000;
	mem[175] = 4'b0000;
	mem[176] = 4'b0000;
	mem[177] = 4'b0000;
	mem[178] = 4'b0000;
	mem[179] = 4'b0000;
	mem[180] = 4'b0000;
	mem[181] = 4'b0000;
	mem[182] = 4'b0000;
	mem[183] = 4'b0000;
	mem[184] = 4'b0000;
	mem[185] = 4'b0000;
	mem[186] = 4'b0000;
	mem[187] = 4'b0000;
	mem[188] = 4'b0000;
	mem[189] = 4'b0000;
	mem[190] = 4'b0000;
	mem[191] = 4'b0000;
	mem[192] = 4'b0000;
	mem[193] = 4'b0000;
	mem[194] = 4'b0000;
	mem[195] = 4'b0000;
	mem[196] = 4'b0000;
	mem[197] = 4'b0000;
	mem[198] = 4'b0000;
	mem[199] = 4'b0000;
	mem[200] = 4'b0000;
	mem[201] = 4'b0000;
	mem[202] = 4'b0000;
	mem[203] = 4'b0000;
	mem[204] = 4'b0000;
	mem[205] = 4'b0000;
	mem[206] = 4'b0000;
	mem[207] = 4'b0000;
	mem[208] = 4'b0000;
	mem[209] = 4'b0000;
	mem[210] = 4'b0000;
	mem[211] = 4'b0000;
	mem[212] = 4'b0000;
	mem[213] = 4'b0000;
	mem[214] = 4'b0000;
	mem[215] = 4'b0000;
	mem[216] = 4'b0000;
	mem[217] = 4'b0000;
	mem[218] = 4'b0000;
	mem[219] = 4'b0000;
	mem[220] = 4'b0000;
	mem[221] = 4'b0000;
	mem[222] = 4'b0000;
	mem[223] = 4'b0000;
	mem[224] = 4'b0000;
	mem[225] = 4'b0000;
	mem[226] = 4'b0000;
	mem[227] = 4'b0000;
	mem[228] = 4'b0000;
	mem[229] = 4'b0000;
	mem[230] = 4'b0000;
	mem[231] = 4'b0000;
	mem[232] = 4'b0000;
	mem[233] = 4'b0000;
	mem[234] = 4'b0000;
	mem[235] = 4'b0000;
	mem[236] = 4'b0000;
	mem[237] = 4'b0000;
	mem[238] = 4'b0000;
	mem[239] = 4'b0000;
	mem[240] = 4'b0000;
	mem[241] = 4'b0000;
	mem[242] = 4'b0000;
	mem[243] = 4'b0000;
	mem[244] = 4'b0000;
	mem[245] = 4'b0000;
	mem[246] = 4'b0000;
	mem[247] = 4'b0000;
	mem[248] = 4'b0000;
	mem[249] = 4'b0000;
	mem[250] = 4'b0000;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0000;
	mem[260] = 4'b0000;
	mem[261] = 4'b0000;
	mem[262] = 4'b0000;
	mem[263] = 4'b0000;
	mem[264] = 4'b0000;
	mem[265] = 4'b0000;
	mem[266] = 4'b0000;
	mem[267] = 4'b0000;
	mem[268] = 4'b0000;
	mem[269] = 4'b0000;
	mem[270] = 4'b0000;
	mem[271] = 4'b0000;
	mem[272] = 4'b0000;
	mem[273] = 4'b0000;
	mem[274] = 4'b0000;
	mem[275] = 4'b0000;
	mem[276] = 4'b0000;
	mem[277] = 4'b0000;
	mem[278] = 4'b0000;
	mem[279] = 4'b0000;
	mem[280] = 4'b0000;
	mem[281] = 4'b0000;
	mem[282] = 4'b0000;
	mem[283] = 4'b0000;
	mem[284] = 4'b0000;
	mem[285] = 4'b0000;
	mem[286] = 4'b0000;
	mem[287] = 4'b0000;
	mem[288] = 4'b0000;
	mem[289] = 4'b0000;
	mem[290] = 4'b0000;
	mem[291] = 4'b0000;
	mem[292] = 4'b0000;
	mem[293] = 4'b0000;
	mem[294] = 4'b0000;
	mem[295] = 4'b0000;
	mem[296] = 4'b0000;
	mem[297] = 4'b0000;
	mem[298] = 4'b0000;
	mem[299] = 4'b0000;
	mem[300] = 4'b0000;
	mem[301] = 4'b0000;
	mem[302] = 4'b0000;
	mem[303] = 4'b0000;
	mem[304] = 4'b0000;
	mem[305] = 4'b0000;
	mem[306] = 4'b0000;
	mem[307] = 4'b0000;
	mem[308] = 4'b0000;
	mem[309] = 4'b0000;
	mem[310] = 4'b0000;
	mem[311] = 4'b0000;
	mem[312] = 4'b0000;
	mem[313] = 4'b0000;
	mem[314] = 4'b0000;
	mem[315] = 4'b0000;
	mem[316] = 4'b0000;
	mem[317] = 4'b0000;
	mem[318] = 4'b0000;
	mem[319] = 4'b0000;
	mem[320] = 4'b0000;
	mem[321] = 4'b0000;
	mem[322] = 4'b0000;
	mem[323] = 4'b0000;
	mem[324] = 4'b0000;
	mem[325] = 4'b0000;
	mem[326] = 4'b0000;
	mem[327] = 4'b0000;
	mem[328] = 4'b0000;
	mem[329] = 4'b0000;
	mem[330] = 4'b0000;
	mem[331] = 4'b0000;
	mem[332] = 4'b0000;
	mem[333] = 4'b0000;
	mem[334] = 4'b0000;
	mem[335] = 4'b0000;
	mem[336] = 4'b0000;
	mem[337] = 4'b0000;
	mem[338] = 4'b0000;
	mem[339] = 4'b0000;
	mem[340] = 4'b0000;
	mem[341] = 4'b0000;
	mem[342] = 4'b0000;
	mem[343] = 4'b0000;
	mem[344] = 4'b0000;
	mem[345] = 4'b0000;
	mem[346] = 4'b0000;
	mem[347] = 4'b0000;
	mem[348] = 4'b0000;
	mem[349] = 4'b0000;
	mem[350] = 4'b0000;
	mem[351] = 4'b0000;
	mem[352] = 4'b0000;
	mem[353] = 4'b0000;
	mem[354] = 4'b0000;
	mem[355] = 4'b0000;
	mem[356] = 4'b0000;
	mem[357] = 4'b0000;
	mem[358] = 4'b0000;
	mem[359] = 4'b0000;
	mem[360] = 4'b0000;
	mem[361] = 4'b0000;
	mem[362] = 4'b0000;
	mem[363] = 4'b0000;
	mem[364] = 4'b0000;
	mem[365] = 4'b0000;
	mem[366] = 4'b0000;
	mem[367] = 4'b0000;
	mem[368] = 4'b0000;
	mem[369] = 4'b0000;
	mem[370] = 4'b0000;
	mem[371] = 4'b0000;
	mem[372] = 4'b0000;
	mem[373] = 4'b0000;
	mem[374] = 4'b0000;
	mem[375] = 4'b0000;
	mem[376] = 4'b0000;
	mem[377] = 4'b0000;
	mem[378] = 4'b0000;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0000;
	mem[388] = 4'b0000;
	mem[389] = 4'b0000;
	mem[390] = 4'b0000;
	mem[391] = 4'b0000;
	mem[392] = 4'b0000;
	mem[393] = 4'b0000;
	mem[394] = 4'b0000;
	mem[395] = 4'b0000;
	mem[396] = 4'b0000;
	mem[397] = 4'b0000;
	mem[398] = 4'b0000;
	mem[399] = 4'b0000;
	mem[400] = 4'b0000;
	mem[401] = 4'b0000;
	mem[402] = 4'b0000;
	mem[403] = 4'b0000;
	mem[404] = 4'b0000;
	mem[405] = 4'b0000;
	mem[406] = 4'b0000;
	mem[407] = 4'b0000;
	mem[408] = 4'b0000;
	mem[409] = 4'b0000;
	mem[410] = 4'b0000;
	mem[411] = 4'b0000;
	mem[412] = 4'b0000;
	mem[413] = 4'b0000;
	mem[414] = 4'b0000;
	mem[415] = 4'b0000;
	mem[416] = 4'b0000;
	mem[417] = 4'b0000;
	mem[418] = 4'b0000;
	mem[419] = 4'b0000;
	mem[420] = 4'b0000;
	mem[421] = 4'b0000;
	mem[422] = 4'b0000;
	mem[423] = 4'b0000;
	mem[424] = 4'b0000;
	mem[425] = 4'b0000;
	mem[426] = 4'b0000;
	mem[427] = 4'b0000;
	mem[428] = 4'b0000;
	mem[429] = 4'b0000;
	mem[430] = 4'b0000;
	mem[431] = 4'b0000;
	mem[432] = 4'b0000;
	mem[433] = 4'b0000;
	mem[434] = 4'b0000;
	mem[435] = 4'b0000;
	mem[436] = 4'b0000;
	mem[437] = 4'b0000;
	mem[438] = 4'b0000;
	mem[439] = 4'b0000;
	mem[440] = 4'b0000;
	mem[441] = 4'b0000;
	mem[442] = 4'b0000;
	mem[443] = 4'b0000;
	mem[444] = 4'b0000;
	mem[445] = 4'b0000;
	mem[446] = 4'b0000;
	mem[447] = 4'b0000;
	mem[448] = 4'b0000;
	mem[449] = 4'b0000;
	mem[450] = 4'b0000;
	mem[451] = 4'b0000;
	mem[452] = 4'b0000;
	mem[453] = 4'b0000;
	mem[454] = 4'b0000;
	mem[455] = 4'b0000;
	mem[456] = 4'b0000;
	mem[457] = 4'b0000;
	mem[458] = 4'b0000;
	mem[459] = 4'b0000;
	mem[460] = 4'b0000;
	mem[461] = 4'b0000;
	mem[462] = 4'b0000;
	mem[463] = 4'b0000;
	mem[464] = 4'b0000;
	mem[465] = 4'b0000;
	mem[466] = 4'b0000;
	mem[467] = 4'b0000;
	mem[468] = 4'b0000;
	mem[469] = 4'b0000;
	mem[470] = 4'b0000;
	mem[471] = 4'b0000;
	mem[472] = 4'b0000;
	mem[473] = 4'b0000;
	mem[474] = 4'b0000;
	mem[475] = 4'b0000;
	mem[476] = 4'b0000;
	mem[477] = 4'b0000;
	mem[478] = 4'b0000;
	mem[479] = 4'b0000;
	mem[480] = 4'b0000;
	mem[481] = 4'b0000;
	mem[482] = 4'b0000;
	mem[483] = 4'b0000;
	mem[484] = 4'b0000;
	mem[485] = 4'b0000;
	mem[486] = 4'b0000;
	mem[487] = 4'b0000;
	mem[488] = 4'b0000;
	mem[489] = 4'b0000;
	mem[490] = 4'b0000;
	mem[491] = 4'b0000;
	mem[492] = 4'b0000;
	mem[493] = 4'b0000;
	mem[494] = 4'b0000;
	mem[495] = 4'b0000;
	mem[496] = 4'b0000;
	mem[497] = 4'b0000;
	mem[498] = 4'b0000;
	mem[499] = 4'b0000;
	mem[500] = 4'b0000;
	mem[501] = 4'b0000;
	mem[502] = 4'b0000;
	mem[503] = 4'b0000;
	mem[504] = 4'b0000;
	mem[505] = 4'b0000;
	mem[506] = 4'b0000;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0000;
	mem[516] = 4'b0000;
	mem[517] = 4'b0000;
	mem[518] = 4'b0000;
	mem[519] = 4'b0000;
	mem[520] = 4'b0000;
	mem[521] = 4'b0000;
	mem[522] = 4'b0000;
	mem[523] = 4'b0000;
	mem[524] = 4'b0000;
	mem[525] = 4'b0000;
	mem[526] = 4'b0000;
	mem[527] = 4'b0000;
	mem[528] = 4'b0000;
	mem[529] = 4'b0000;
	mem[530] = 4'b0000;
	mem[531] = 4'b0000;
	mem[532] = 4'b0000;
	mem[533] = 4'b0000;
	mem[534] = 4'b0000;
	mem[535] = 4'b0000;
	mem[536] = 4'b0000;
	mem[537] = 4'b0000;
	mem[538] = 4'b0000;
	mem[539] = 4'b0000;
	mem[540] = 4'b0000;
	mem[541] = 4'b0000;
	mem[542] = 4'b0000;
	mem[543] = 4'b0000;
	mem[544] = 4'b0000;
	mem[545] = 4'b0000;
	mem[546] = 4'b0000;
	mem[547] = 4'b0000;
	mem[548] = 4'b0000;
	mem[549] = 4'b0000;
	mem[550] = 4'b0000;
	mem[551] = 4'b0000;
	mem[552] = 4'b0000;
	mem[553] = 4'b0000;
	mem[554] = 4'b0000;
	mem[555] = 4'b0000;
	mem[556] = 4'b0000;
	mem[557] = 4'b0000;
	mem[558] = 4'b0000;
	mem[559] = 4'b0000;
	mem[560] = 4'b0000;
	mem[561] = 4'b0000;
	mem[562] = 4'b0000;
	mem[563] = 4'b0000;
	mem[564] = 4'b0000;
	mem[565] = 4'b0000;
	mem[566] = 4'b0000;
	mem[567] = 4'b0000;
	mem[568] = 4'b0000;
	mem[569] = 4'b0000;
	mem[570] = 4'b0000;
	mem[571] = 4'b0000;
	mem[572] = 4'b0000;
	mem[573] = 4'b0000;
	mem[574] = 4'b0000;
	mem[575] = 4'b0000;
	mem[576] = 4'b0000;
	mem[577] = 4'b0000;
	mem[578] = 4'b0000;
	mem[579] = 4'b0000;
	mem[580] = 4'b0000;
	mem[581] = 4'b0000;
	mem[582] = 4'b0000;
	mem[583] = 4'b0000;
	mem[584] = 4'b0000;
	mem[585] = 4'b0000;
	mem[586] = 4'b0000;
	mem[587] = 4'b0000;
	mem[588] = 4'b0000;
	mem[589] = 4'b0000;
	mem[590] = 4'b0000;
	mem[591] = 4'b0000;
	mem[592] = 4'b0000;
	mem[593] = 4'b0000;
	mem[594] = 4'b0000;
	mem[595] = 4'b0000;
	mem[596] = 4'b0000;
	mem[597] = 4'b0000;
	mem[598] = 4'b0000;
	mem[599] = 4'b0000;
	mem[600] = 4'b0000;
	mem[601] = 4'b0000;
	mem[602] = 4'b0000;
	mem[603] = 4'b0000;
	mem[604] = 4'b0000;
	mem[605] = 4'b0000;
	mem[606] = 4'b0000;
	mem[607] = 4'b0000;
	mem[608] = 4'b0000;
	mem[609] = 4'b0000;
	mem[610] = 4'b0000;
	mem[611] = 4'b0000;
	mem[612] = 4'b0000;
	mem[613] = 4'b0000;
	mem[614] = 4'b0000;
	mem[615] = 4'b0000;
	mem[616] = 4'b0000;
	mem[617] = 4'b0000;
	mem[618] = 4'b0000;
	mem[619] = 4'b0000;
	mem[620] = 4'b0000;
	mem[621] = 4'b0000;
	mem[622] = 4'b0000;
	mem[623] = 4'b0000;
	mem[624] = 4'b0000;
	mem[625] = 4'b0000;
	mem[626] = 4'b0000;
	mem[627] = 4'b0000;
	mem[628] = 4'b0000;
	mem[629] = 4'b0000;
	mem[630] = 4'b0000;
	mem[631] = 4'b0000;
	mem[632] = 4'b0000;
	mem[633] = 4'b0000;
	mem[634] = 4'b0000;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0000;
	mem[644] = 4'b0000;
	mem[645] = 4'b0000;
	mem[646] = 4'b0000;
	mem[647] = 4'b0000;
	mem[648] = 4'b0000;
	mem[649] = 4'b0000;
	mem[650] = 4'b0000;
	mem[651] = 4'b0000;
	mem[652] = 4'b0000;
	mem[653] = 4'b0000;
	mem[654] = 4'b0000;
	mem[655] = 4'b0000;
	mem[656] = 4'b0000;
	mem[657] = 4'b0000;
	mem[658] = 4'b0000;
	mem[659] = 4'b0000;
	mem[660] = 4'b0000;
	mem[661] = 4'b0000;
	mem[662] = 4'b0000;
	mem[663] = 4'b0000;
	mem[664] = 4'b0000;
	mem[665] = 4'b0000;
	mem[666] = 4'b0000;
	mem[667] = 4'b0000;
	mem[668] = 4'b0000;
	mem[669] = 4'b0000;
	mem[670] = 4'b0000;
	mem[671] = 4'b0000;
	mem[672] = 4'b0000;
	mem[673] = 4'b0000;
	mem[674] = 4'b0000;
	mem[675] = 4'b0000;
	mem[676] = 4'b0000;
	mem[677] = 4'b0000;
	mem[678] = 4'b0000;
	mem[679] = 4'b0000;
	mem[680] = 4'b0000;
	mem[681] = 4'b0000;
	mem[682] = 4'b0000;
	mem[683] = 4'b0000;
	mem[684] = 4'b0000;
	mem[685] = 4'b0000;
	mem[686] = 4'b0000;
	mem[687] = 4'b0000;
	mem[688] = 4'b0000;
	mem[689] = 4'b0000;
	mem[690] = 4'b0000;
	mem[691] = 4'b0000;
	mem[692] = 4'b0000;
	mem[693] = 4'b0000;
	mem[694] = 4'b0000;
	mem[695] = 4'b0000;
	mem[696] = 4'b0000;
	mem[697] = 4'b0000;
	mem[698] = 4'b0000;
	mem[699] = 4'b0000;
	mem[700] = 4'b0000;
	mem[701] = 4'b0000;
	mem[702] = 4'b0000;
	mem[703] = 4'b0000;
	mem[704] = 4'b0000;
	mem[705] = 4'b0000;
	mem[706] = 4'b0000;
	mem[707] = 4'b0000;
	mem[708] = 4'b0000;
	mem[709] = 4'b0000;
	mem[710] = 4'b0000;
	mem[711] = 4'b0000;
	mem[712] = 4'b0000;
	mem[713] = 4'b0000;
	mem[714] = 4'b0000;
	mem[715] = 4'b0000;
	mem[716] = 4'b0000;
	mem[717] = 4'b0000;
	mem[718] = 4'b0000;
	mem[719] = 4'b0000;
	mem[720] = 4'b0000;
	mem[721] = 4'b0000;
	mem[722] = 4'b0000;
	mem[723] = 4'b0000;
	mem[724] = 4'b0000;
	mem[725] = 4'b0000;
	mem[726] = 4'b0000;
	mem[727] = 4'b0000;
	mem[728] = 4'b0000;
	mem[729] = 4'b0000;
	mem[730] = 4'b0000;
	mem[731] = 4'b0000;
	mem[732] = 4'b0000;
	mem[733] = 4'b0000;
	mem[734] = 4'b0000;
	mem[735] = 4'b0000;
	mem[736] = 4'b0000;
	mem[737] = 4'b0000;
	mem[738] = 4'b0000;
	mem[739] = 4'b0000;
	mem[740] = 4'b0000;
	mem[741] = 4'b0000;
	mem[742] = 4'b0000;
	mem[743] = 4'b0000;
	mem[744] = 4'b0000;
	mem[745] = 4'b0000;
	mem[746] = 4'b0000;
	mem[747] = 4'b0000;
	mem[748] = 4'b0000;
	mem[749] = 4'b0000;
	mem[750] = 4'b0000;
	mem[751] = 4'b0000;
	mem[752] = 4'b0000;
	mem[753] = 4'b0000;
	mem[754] = 4'b0000;
	mem[755] = 4'b0000;
	mem[756] = 4'b0000;
	mem[757] = 4'b0000;
	mem[758] = 4'b0000;
	mem[759] = 4'b0000;
	mem[760] = 4'b0000;
	mem[761] = 4'b0000;
	mem[762] = 4'b0000;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0000;
	mem[772] = 4'b0000;
	mem[773] = 4'b0000;
	mem[774] = 4'b0000;
	mem[775] = 4'b0000;
	mem[776] = 4'b0000;
	mem[777] = 4'b0000;
	mem[778] = 4'b0000;
	mem[779] = 4'b0000;
	mem[780] = 4'b0000;
	mem[781] = 4'b0000;
	mem[782] = 4'b0000;
	mem[783] = 4'b0000;
	mem[784] = 4'b0000;
	mem[785] = 4'b0000;
	mem[786] = 4'b0000;
	mem[787] = 4'b0000;
	mem[788] = 4'b0000;
	mem[789] = 4'b0000;
	mem[790] = 4'b0000;
	mem[791] = 4'b0000;
	mem[792] = 4'b0000;
	mem[793] = 4'b0000;
	mem[794] = 4'b0000;
	mem[795] = 4'b0000;
	mem[796] = 4'b0000;
	mem[797] = 4'b0000;
	mem[798] = 4'b0000;
	mem[799] = 4'b0000;
	mem[800] = 4'b0000;
	mem[801] = 4'b0000;
	mem[802] = 4'b0000;
	mem[803] = 4'b0000;
	mem[804] = 4'b0000;
	mem[805] = 4'b0000;
	mem[806] = 4'b0000;
	mem[807] = 4'b0000;
	mem[808] = 4'b0000;
	mem[809] = 4'b0000;
	mem[810] = 4'b0000;
	mem[811] = 4'b0000;
	mem[812] = 4'b0000;
	mem[813] = 4'b0000;
	mem[814] = 4'b0000;
	mem[815] = 4'b0000;
	mem[816] = 4'b0000;
	mem[817] = 4'b0000;
	mem[818] = 4'b0000;
	mem[819] = 4'b0000;
	mem[820] = 4'b0000;
	mem[821] = 4'b0000;
	mem[822] = 4'b0000;
	mem[823] = 4'b0000;
	mem[824] = 4'b0000;
	mem[825] = 4'b0000;
	mem[826] = 4'b0000;
	mem[827] = 4'b0000;
	mem[828] = 4'b0000;
	mem[829] = 4'b0000;
	mem[830] = 4'b0000;
	mem[831] = 4'b0000;
	mem[832] = 4'b0000;
	mem[833] = 4'b0000;
	mem[834] = 4'b0000;
	mem[835] = 4'b0000;
	mem[836] = 4'b0000;
	mem[837] = 4'b0000;
	mem[838] = 4'b0000;
	mem[839] = 4'b0000;
	mem[840] = 4'b0000;
	mem[841] = 4'b0000;
	mem[842] = 4'b0000;
	mem[843] = 4'b0000;
	mem[844] = 4'b0000;
	mem[845] = 4'b0000;
	mem[846] = 4'b0000;
	mem[847] = 4'b0000;
	mem[848] = 4'b0000;
	mem[849] = 4'b0000;
	mem[850] = 4'b0000;
	mem[851] = 4'b0000;
	mem[852] = 4'b0000;
	mem[853] = 4'b0000;
	mem[854] = 4'b0000;
	mem[855] = 4'b0000;
	mem[856] = 4'b0000;
	mem[857] = 4'b0000;
	mem[858] = 4'b0000;
	mem[859] = 4'b0000;
	mem[860] = 4'b0000;
	mem[861] = 4'b0000;
	mem[862] = 4'b0000;
	mem[863] = 4'b0000;
	mem[864] = 4'b0000;
	mem[865] = 4'b0000;
	mem[866] = 4'b0000;
	mem[867] = 4'b0000;
	mem[868] = 4'b0000;
	mem[869] = 4'b0000;
	mem[870] = 4'b0000;
	mem[871] = 4'b0000;
	mem[872] = 4'b0000;
	mem[873] = 4'b0000;
	mem[874] = 4'b0000;
	mem[875] = 4'b0000;
	mem[876] = 4'b0000;
	mem[877] = 4'b0000;
	mem[878] = 4'b0000;
	mem[879] = 4'b0000;
	mem[880] = 4'b0000;
	mem[881] = 4'b0000;
	mem[882] = 4'b0000;
	mem[883] = 4'b0000;
	mem[884] = 4'b0000;
	mem[885] = 4'b0000;
	mem[886] = 4'b0000;
	mem[887] = 4'b0000;
	mem[888] = 4'b0000;
	mem[889] = 4'b0000;
	mem[890] = 4'b0000;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0000;
	mem[900] = 4'b0000;
	mem[901] = 4'b0000;
	mem[902] = 4'b0000;
	mem[903] = 4'b0000;
	mem[904] = 4'b0000;
	mem[905] = 4'b0000;
	mem[906] = 4'b0000;
	mem[907] = 4'b0000;
	mem[908] = 4'b0000;
	mem[909] = 4'b0000;
	mem[910] = 4'b0000;
	mem[911] = 4'b0000;
	mem[912] = 4'b0000;
	mem[913] = 4'b0000;
	mem[914] = 4'b0000;
	mem[915] = 4'b0000;
	mem[916] = 4'b0000;
	mem[917] = 4'b0000;
	mem[918] = 4'b0000;
	mem[919] = 4'b0000;
	mem[920] = 4'b0000;
	mem[921] = 4'b0000;
	mem[922] = 4'b0000;
	mem[923] = 4'b0000;
	mem[924] = 4'b0000;
	mem[925] = 4'b0000;
	mem[926] = 4'b0000;
	mem[927] = 4'b0000;
	mem[928] = 4'b0000;
	mem[929] = 4'b0000;
	mem[930] = 4'b0000;
	mem[931] = 4'b0000;
	mem[932] = 4'b0000;
	mem[933] = 4'b0000;
	mem[934] = 4'b0000;
	mem[935] = 4'b0000;
	mem[936] = 4'b0000;
	mem[937] = 4'b0000;
	mem[938] = 4'b0000;
	mem[939] = 4'b0000;
	mem[940] = 4'b0000;
	mem[941] = 4'b0000;
	mem[942] = 4'b0000;
	mem[943] = 4'b0000;
	mem[944] = 4'b0000;
	mem[945] = 4'b0000;
	mem[946] = 4'b0000;
	mem[947] = 4'b0000;
	mem[948] = 4'b0000;
	mem[949] = 4'b0000;
	mem[950] = 4'b0000;
	mem[951] = 4'b0000;
	mem[952] = 4'b0000;
	mem[953] = 4'b0000;
	mem[954] = 4'b0000;
	mem[955] = 4'b0000;
	mem[956] = 4'b0000;
	mem[957] = 4'b0000;
	mem[958] = 4'b0000;
	mem[959] = 4'b0000;
	mem[960] = 4'b0000;
	mem[961] = 4'b0000;
	mem[962] = 4'b0000;
	mem[963] = 4'b0000;
	mem[964] = 4'b0000;
	mem[965] = 4'b0000;
	mem[966] = 4'b0000;
	mem[967] = 4'b0000;
	mem[968] = 4'b0000;
	mem[969] = 4'b0000;
	mem[970] = 4'b0000;
	mem[971] = 4'b0000;
	mem[972] = 4'b0000;
	mem[973] = 4'b0000;
	mem[974] = 4'b0000;
	mem[975] = 4'b0000;
	mem[976] = 4'b0000;
	mem[977] = 4'b0000;
	mem[978] = 4'b0000;
	mem[979] = 4'b0000;
	mem[980] = 4'b0000;
	mem[981] = 4'b0000;
	mem[982] = 4'b0000;
	mem[983] = 4'b0000;
	mem[984] = 4'b0000;
	mem[985] = 4'b0000;
	mem[986] = 4'b0000;
	mem[987] = 4'b0000;
	mem[988] = 4'b0000;
	mem[989] = 4'b0000;
	mem[990] = 4'b0000;
	mem[991] = 4'b0000;
	mem[992] = 4'b0000;
	mem[993] = 4'b0000;
	mem[994] = 4'b0000;
	mem[995] = 4'b0000;
	mem[996] = 4'b0000;
	mem[997] = 4'b0000;
	mem[998] = 4'b0000;
	mem[999] = 4'b0000;
	mem[1000] = 4'b0000;
	mem[1001] = 4'b0000;
	mem[1002] = 4'b0000;
	mem[1003] = 4'b0000;
	mem[1004] = 4'b0000;
	mem[1005] = 4'b0000;
	mem[1006] = 4'b0000;
	mem[1007] = 4'b0000;
	mem[1008] = 4'b0000;
	mem[1009] = 4'b0000;
	mem[1010] = 4'b0000;
	mem[1011] = 4'b0000;
	mem[1012] = 4'b0000;
	mem[1013] = 4'b0000;
	mem[1014] = 4'b0000;
	mem[1015] = 4'b0000;
	mem[1016] = 4'b0000;
	mem[1017] = 4'b0000;
	mem[1018] = 4'b0000;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0000;
	mem[1028] = 4'b0000;
	mem[1029] = 4'b0000;
	mem[1030] = 4'b0000;
	mem[1031] = 4'b0000;
	mem[1032] = 4'b0000;
	mem[1033] = 4'b0000;
	mem[1034] = 4'b0000;
	mem[1035] = 4'b0000;
	mem[1036] = 4'b0000;
	mem[1037] = 4'b0000;
	mem[1038] = 4'b0000;
	mem[1039] = 4'b0000;
	mem[1040] = 4'b0000;
	mem[1041] = 4'b0000;
	mem[1042] = 4'b0000;
	mem[1043] = 4'b0000;
	mem[1044] = 4'b0000;
	mem[1045] = 4'b0000;
	mem[1046] = 4'b0000;
	mem[1047] = 4'b0000;
	mem[1048] = 4'b0000;
	mem[1049] = 4'b0000;
	mem[1050] = 4'b0000;
	mem[1051] = 4'b0000;
	mem[1052] = 4'b0000;
	mem[1053] = 4'b0000;
	mem[1054] = 4'b0000;
	mem[1055] = 4'b0000;
	mem[1056] = 4'b0000;
	mem[1057] = 4'b0000;
	mem[1058] = 4'b0000;
	mem[1059] = 4'b0000;
	mem[1060] = 4'b0000;
	mem[1061] = 4'b0000;
	mem[1062] = 4'b0000;
	mem[1063] = 4'b0000;
	mem[1064] = 4'b0000;
	mem[1065] = 4'b0000;
	mem[1066] = 4'b0000;
	mem[1067] = 4'b0000;
	mem[1068] = 4'b0000;
	mem[1069] = 4'b0000;
	mem[1070] = 4'b0000;
	mem[1071] = 4'b0000;
	mem[1072] = 4'b0000;
	mem[1073] = 4'b0000;
	mem[1074] = 4'b0000;
	mem[1075] = 4'b0000;
	mem[1076] = 4'b0000;
	mem[1077] = 4'b0000;
	mem[1078] = 4'b0000;
	mem[1079] = 4'b0000;
	mem[1080] = 4'b0000;
	mem[1081] = 4'b0000;
	mem[1082] = 4'b0000;
	mem[1083] = 4'b0000;
	mem[1084] = 4'b0000;
	mem[1085] = 4'b0000;
	mem[1086] = 4'b0000;
	mem[1087] = 4'b0000;
	mem[1088] = 4'b0000;
	mem[1089] = 4'b0001;
	mem[1090] = 4'b0001;
	mem[1091] = 4'b0000;
	mem[1092] = 4'b0000;
	mem[1093] = 4'b0000;
	mem[1094] = 4'b0000;
	mem[1095] = 4'b0000;
	mem[1096] = 4'b0000;
	mem[1097] = 4'b0000;
	mem[1098] = 4'b0000;
	mem[1099] = 4'b0000;
	mem[1100] = 4'b0000;
	mem[1101] = 4'b0000;
	mem[1102] = 4'b0000;
	mem[1103] = 4'b0000;
	mem[1104] = 4'b0000;
	mem[1105] = 4'b0000;
	mem[1106] = 4'b0000;
	mem[1107] = 4'b0000;
	mem[1108] = 4'b0000;
	mem[1109] = 4'b0000;
	mem[1110] = 4'b0000;
	mem[1111] = 4'b0000;
	mem[1112] = 4'b0000;
	mem[1113] = 4'b0000;
	mem[1114] = 4'b0000;
	mem[1115] = 4'b0000;
	mem[1116] = 4'b0000;
	mem[1117] = 4'b0000;
	mem[1118] = 4'b0000;
	mem[1119] = 4'b0000;
	mem[1120] = 4'b0000;
	mem[1121] = 4'b0000;
	mem[1122] = 4'b0000;
	mem[1123] = 4'b0000;
	mem[1124] = 4'b0000;
	mem[1125] = 4'b0000;
	mem[1126] = 4'b0000;
	mem[1127] = 4'b0000;
	mem[1128] = 4'b0000;
	mem[1129] = 4'b0000;
	mem[1130] = 4'b0000;
	mem[1131] = 4'b0000;
	mem[1132] = 4'b0000;
	mem[1133] = 4'b0000;
	mem[1134] = 4'b0000;
	mem[1135] = 4'b0000;
	mem[1136] = 4'b0000;
	mem[1137] = 4'b0000;
	mem[1138] = 4'b0000;
	mem[1139] = 4'b0000;
	mem[1140] = 4'b0000;
	mem[1141] = 4'b0000;
	mem[1142] = 4'b0000;
	mem[1143] = 4'b0000;
	mem[1144] = 4'b0000;
	mem[1145] = 4'b0000;
	mem[1146] = 4'b0000;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0000;
	mem[1156] = 4'b0000;
	mem[1157] = 4'b0000;
	mem[1158] = 4'b0000;
	mem[1159] = 4'b0000;
	mem[1160] = 4'b0000;
	mem[1161] = 4'b0000;
	mem[1162] = 4'b0000;
	mem[1163] = 4'b0000;
	mem[1164] = 4'b0000;
	mem[1165] = 4'b0000;
	mem[1166] = 4'b0000;
	mem[1167] = 4'b0000;
	mem[1168] = 4'b0000;
	mem[1169] = 4'b0000;
	mem[1170] = 4'b0000;
	mem[1171] = 4'b0000;
	mem[1172] = 4'b0000;
	mem[1173] = 4'b0000;
	mem[1174] = 4'b0000;
	mem[1175] = 4'b0000;
	mem[1176] = 4'b0000;
	mem[1177] = 4'b0000;
	mem[1178] = 4'b0000;
	mem[1179] = 4'b0000;
	mem[1180] = 4'b0000;
	mem[1181] = 4'b0000;
	mem[1182] = 4'b0000;
	mem[1183] = 4'b0000;
	mem[1184] = 4'b0000;
	mem[1185] = 4'b0000;
	mem[1186] = 4'b0000;
	mem[1187] = 4'b0000;
	mem[1188] = 4'b0000;
	mem[1189] = 4'b0000;
	mem[1190] = 4'b0000;
	mem[1191] = 4'b0000;
	mem[1192] = 4'b0000;
	mem[1193] = 4'b0000;
	mem[1194] = 4'b0000;
	mem[1195] = 4'b0000;
	mem[1196] = 4'b0000;
	mem[1197] = 4'b0000;
	mem[1198] = 4'b0000;
	mem[1199] = 4'b0000;
	mem[1200] = 4'b0000;
	mem[1201] = 4'b0000;
	mem[1202] = 4'b0000;
	mem[1203] = 4'b0000;
	mem[1204] = 4'b0000;
	mem[1205] = 4'b0000;
	mem[1206] = 4'b0000;
	mem[1207] = 4'b0000;
	mem[1208] = 4'b0000;
	mem[1209] = 4'b0000;
	mem[1210] = 4'b0000;
	mem[1211] = 4'b0000;
	mem[1212] = 4'b0000;
	mem[1213] = 4'b0000;
	mem[1214] = 4'b0000;
	mem[1215] = 4'b0000;
	mem[1216] = 4'b0001;
	mem[1217] = 4'b0001;
	mem[1218] = 4'b0000;
	mem[1219] = 4'b0000;
	mem[1220] = 4'b0000;
	mem[1221] = 4'b0000;
	mem[1222] = 4'b0000;
	mem[1223] = 4'b0000;
	mem[1224] = 4'b0000;
	mem[1225] = 4'b0000;
	mem[1226] = 4'b0000;
	mem[1227] = 4'b0000;
	mem[1228] = 4'b0000;
	mem[1229] = 4'b0000;
	mem[1230] = 4'b0000;
	mem[1231] = 4'b0000;
	mem[1232] = 4'b0000;
	mem[1233] = 4'b0000;
	mem[1234] = 4'b0000;
	mem[1235] = 4'b0000;
	mem[1236] = 4'b0000;
	mem[1237] = 4'b0000;
	mem[1238] = 4'b0000;
	mem[1239] = 4'b0000;
	mem[1240] = 4'b0000;
	mem[1241] = 4'b0000;
	mem[1242] = 4'b0000;
	mem[1243] = 4'b0000;
	mem[1244] = 4'b0000;
	mem[1245] = 4'b0000;
	mem[1246] = 4'b0000;
	mem[1247] = 4'b0000;
	mem[1248] = 4'b0000;
	mem[1249] = 4'b0000;
	mem[1250] = 4'b0000;
	mem[1251] = 4'b0000;
	mem[1252] = 4'b0000;
	mem[1253] = 4'b0000;
	mem[1254] = 4'b0000;
	mem[1255] = 4'b0000;
	mem[1256] = 4'b0000;
	mem[1257] = 4'b0000;
	mem[1258] = 4'b0000;
	mem[1259] = 4'b0000;
	mem[1260] = 4'b0000;
	mem[1261] = 4'b0000;
	mem[1262] = 4'b0000;
	mem[1263] = 4'b0000;
	mem[1264] = 4'b0000;
	mem[1265] = 4'b0000;
	mem[1266] = 4'b0000;
	mem[1267] = 4'b0000;
	mem[1268] = 4'b0000;
	mem[1269] = 4'b0000;
	mem[1270] = 4'b0000;
	mem[1271] = 4'b0000;
	mem[1272] = 4'b0000;
	mem[1273] = 4'b0000;
	mem[1274] = 4'b0000;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0000;
	mem[1284] = 4'b0000;
	mem[1285] = 4'b0000;
	mem[1286] = 4'b0000;
	mem[1287] = 4'b0000;
	mem[1288] = 4'b0000;
	mem[1289] = 4'b0000;
	mem[1290] = 4'b0000;
	mem[1291] = 4'b0000;
	mem[1292] = 4'b0000;
	mem[1293] = 4'b0000;
	mem[1294] = 4'b0000;
	mem[1295] = 4'b0000;
	mem[1296] = 4'b0000;
	mem[1297] = 4'b0000;
	mem[1298] = 4'b0000;
	mem[1299] = 4'b0000;
	mem[1300] = 4'b0000;
	mem[1301] = 4'b0000;
	mem[1302] = 4'b0000;
	mem[1303] = 4'b0000;
	mem[1304] = 4'b0000;
	mem[1305] = 4'b0000;
	mem[1306] = 4'b0000;
	mem[1307] = 4'b0000;
	mem[1308] = 4'b0000;
	mem[1309] = 4'b0000;
	mem[1310] = 4'b0000;
	mem[1311] = 4'b0000;
	mem[1312] = 4'b0000;
	mem[1313] = 4'b0000;
	mem[1314] = 4'b0000;
	mem[1315] = 4'b0000;
	mem[1316] = 4'b0000;
	mem[1317] = 4'b0000;
	mem[1318] = 4'b0000;
	mem[1319] = 4'b0000;
	mem[1320] = 4'b0000;
	mem[1321] = 4'b0000;
	mem[1322] = 4'b0000;
	mem[1323] = 4'b0000;
	mem[1324] = 4'b0000;
	mem[1325] = 4'b0000;
	mem[1326] = 4'b0000;
	mem[1327] = 4'b0000;
	mem[1328] = 4'b0000;
	mem[1329] = 4'b0000;
	mem[1330] = 4'b0000;
	mem[1331] = 4'b0000;
	mem[1332] = 4'b0000;
	mem[1333] = 4'b0000;
	mem[1334] = 4'b0000;
	mem[1335] = 4'b0000;
	mem[1336] = 4'b0000;
	mem[1337] = 4'b0000;
	mem[1338] = 4'b0000;
	mem[1339] = 4'b0000;
	mem[1340] = 4'b0000;
	mem[1341] = 4'b0000;
	mem[1342] = 4'b0000;
	mem[1343] = 4'b0000;
	mem[1344] = 4'b0001;
	mem[1345] = 4'b0000;
	mem[1346] = 4'b0000;
	mem[1347] = 4'b0000;
	mem[1348] = 4'b0000;
	mem[1349] = 4'b0000;
	mem[1350] = 4'b0000;
	mem[1351] = 4'b0000;
	mem[1352] = 4'b0000;
	mem[1353] = 4'b0000;
	mem[1354] = 4'b0000;
	mem[1355] = 4'b0000;
	mem[1356] = 4'b0000;
	mem[1357] = 4'b0000;
	mem[1358] = 4'b0000;
	mem[1359] = 4'b0000;
	mem[1360] = 4'b0000;
	mem[1361] = 4'b0000;
	mem[1362] = 4'b0000;
	mem[1363] = 4'b0000;
	mem[1364] = 4'b0000;
	mem[1365] = 4'b0000;
	mem[1366] = 4'b0000;
	mem[1367] = 4'b0000;
	mem[1368] = 4'b0000;
	mem[1369] = 4'b0000;
	mem[1370] = 4'b0000;
	mem[1371] = 4'b0000;
	mem[1372] = 4'b0000;
	mem[1373] = 4'b0000;
	mem[1374] = 4'b0000;
	mem[1375] = 4'b0000;
	mem[1376] = 4'b0000;
	mem[1377] = 4'b0000;
	mem[1378] = 4'b0000;
	mem[1379] = 4'b0000;
	mem[1380] = 4'b0000;
	mem[1381] = 4'b0000;
	mem[1382] = 4'b0000;
	mem[1383] = 4'b0000;
	mem[1384] = 4'b0000;
	mem[1385] = 4'b0000;
	mem[1386] = 4'b0000;
	mem[1387] = 4'b0000;
	mem[1388] = 4'b0000;
	mem[1389] = 4'b0000;
	mem[1390] = 4'b0000;
	mem[1391] = 4'b0000;
	mem[1392] = 4'b0000;
	mem[1393] = 4'b0000;
	mem[1394] = 4'b0000;
	mem[1395] = 4'b0000;
	mem[1396] = 4'b0000;
	mem[1397] = 4'b0000;
	mem[1398] = 4'b0000;
	mem[1399] = 4'b0000;
	mem[1400] = 4'b0000;
	mem[1401] = 4'b0000;
	mem[1402] = 4'b0000;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0101;
	mem[1412] = 4'b0111;
	mem[1413] = 4'b0111;
	mem[1414] = 4'b0111;
	mem[1415] = 4'b0111;
	mem[1416] = 4'b0111;
	mem[1417] = 4'b0111;
	mem[1418] = 4'b0111;
	mem[1419] = 4'b0111;
	mem[1420] = 4'b0111;
	mem[1421] = 4'b0111;
	mem[1422] = 4'b0111;
	mem[1423] = 4'b0111;
	mem[1424] = 4'b0111;
	mem[1425] = 4'b0111;
	mem[1426] = 4'b0111;
	mem[1427] = 4'b0111;
	mem[1428] = 4'b1001;
	mem[1429] = 4'b1001;
	mem[1430] = 4'b1001;
	mem[1431] = 4'b1001;
	mem[1432] = 4'b1001;
	mem[1433] = 4'b1001;
	mem[1434] = 4'b1001;
	mem[1435] = 4'b1001;
	mem[1436] = 4'b1001;
	mem[1437] = 4'b1001;
	mem[1438] = 4'b1001;
	mem[1439] = 4'b1001;
	mem[1440] = 4'b1001;
	mem[1441] = 4'b1001;
	mem[1442] = 4'b1001;
	mem[1443] = 4'b1001;
	mem[1444] = 4'b1001;
	mem[1445] = 4'b1001;
	mem[1446] = 4'b1001;
	mem[1447] = 4'b1001;
	mem[1448] = 4'b1001;
	mem[1449] = 4'b1001;
	mem[1450] = 4'b1001;
	mem[1451] = 4'b1001;
	mem[1452] = 4'b1001;
	mem[1453] = 4'b1001;
	mem[1454] = 4'b1001;
	mem[1455] = 4'b1001;
	mem[1456] = 4'b1001;
	mem[1457] = 4'b1001;
	mem[1458] = 4'b1001;
	mem[1459] = 4'b1001;
	mem[1460] = 4'b1001;
	mem[1461] = 4'b1001;
	mem[1462] = 4'b1001;
	mem[1463] = 4'b1001;
	mem[1464] = 4'b1001;
	mem[1465] = 4'b1001;
	mem[1466] = 4'b1001;
	mem[1467] = 4'b1001;
	mem[1468] = 4'b1001;
	mem[1469] = 4'b1001;
	mem[1470] = 4'b1001;
	mem[1471] = 4'b1000;
	mem[1472] = 4'b1001;
	mem[1473] = 4'b1010;
	mem[1474] = 4'b1001;
	mem[1475] = 4'b1001;
	mem[1476] = 4'b1001;
	mem[1477] = 4'b1001;
	mem[1478] = 4'b1000;
	mem[1479] = 4'b0010;
	mem[1480] = 4'b0001;
	mem[1481] = 4'b0000;
	mem[1482] = 4'b0000;
	mem[1483] = 4'b0000;
	mem[1484] = 4'b0000;
	mem[1485] = 4'b0000;
	mem[1486] = 4'b0000;
	mem[1487] = 4'b0000;
	mem[1488] = 4'b0000;
	mem[1489] = 4'b0000;
	mem[1490] = 4'b0000;
	mem[1491] = 4'b0000;
	mem[1492] = 4'b0000;
	mem[1493] = 4'b0000;
	mem[1494] = 4'b0000;
	mem[1495] = 4'b0000;
	mem[1496] = 4'b0000;
	mem[1497] = 4'b0000;
	mem[1498] = 4'b0000;
	mem[1499] = 4'b0000;
	mem[1500] = 4'b0000;
	mem[1501] = 4'b0000;
	mem[1502] = 4'b0000;
	mem[1503] = 4'b0000;
	mem[1504] = 4'b0000;
	mem[1505] = 4'b0000;
	mem[1506] = 4'b0000;
	mem[1507] = 4'b0000;
	mem[1508] = 4'b0000;
	mem[1509] = 4'b0000;
	mem[1510] = 4'b0000;
	mem[1511] = 4'b0000;
	mem[1512] = 4'b0000;
	mem[1513] = 4'b0000;
	mem[1514] = 4'b0000;
	mem[1515] = 4'b0000;
	mem[1516] = 4'b0000;
	mem[1517] = 4'b0000;
	mem[1518] = 4'b0000;
	mem[1519] = 4'b0000;
	mem[1520] = 4'b0000;
	mem[1521] = 4'b0000;
	mem[1522] = 4'b0000;
	mem[1523] = 4'b0000;
	mem[1524] = 4'b0000;
	mem[1525] = 4'b0000;
	mem[1526] = 4'b0000;
	mem[1527] = 4'b0000;
	mem[1528] = 4'b0000;
	mem[1529] = 4'b0000;
	mem[1530] = 4'b0000;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0111;
	mem[1540] = 4'b1100;
	mem[1541] = 4'b1100;
	mem[1542] = 4'b1100;
	mem[1543] = 4'b1100;
	mem[1544] = 4'b1100;
	mem[1545] = 4'b1100;
	mem[1546] = 4'b1100;
	mem[1547] = 4'b1100;
	mem[1548] = 4'b1100;
	mem[1549] = 4'b1100;
	mem[1550] = 4'b1100;
	mem[1551] = 4'b1100;
	mem[1552] = 4'b1100;
	mem[1553] = 4'b1100;
	mem[1554] = 4'b1100;
	mem[1555] = 4'b1100;
	mem[1556] = 4'b1111;
	mem[1557] = 4'b1111;
	mem[1558] = 4'b1111;
	mem[1559] = 4'b1111;
	mem[1560] = 4'b1111;
	mem[1561] = 4'b1111;
	mem[1562] = 4'b1111;
	mem[1563] = 4'b1111;
	mem[1564] = 4'b1111;
	mem[1565] = 4'b1111;
	mem[1566] = 4'b1111;
	mem[1567] = 4'b1111;
	mem[1568] = 4'b1111;
	mem[1569] = 4'b1111;
	mem[1570] = 4'b1111;
	mem[1571] = 4'b1111;
	mem[1572] = 4'b1111;
	mem[1573] = 4'b1111;
	mem[1574] = 4'b1111;
	mem[1575] = 4'b1111;
	mem[1576] = 4'b1111;
	mem[1577] = 4'b1111;
	mem[1578] = 4'b1111;
	mem[1579] = 4'b1111;
	mem[1580] = 4'b1111;
	mem[1581] = 4'b1111;
	mem[1582] = 4'b1111;
	mem[1583] = 4'b1111;
	mem[1584] = 4'b1111;
	mem[1585] = 4'b1111;
	mem[1586] = 4'b1111;
	mem[1587] = 4'b1111;
	mem[1588] = 4'b1111;
	mem[1589] = 4'b1111;
	mem[1590] = 4'b1111;
	mem[1591] = 4'b1111;
	mem[1592] = 4'b1111;
	mem[1593] = 4'b1111;
	mem[1594] = 4'b1111;
	mem[1595] = 4'b1111;
	mem[1596] = 4'b1111;
	mem[1597] = 4'b1111;
	mem[1598] = 4'b1111;
	mem[1599] = 4'b1101;
	mem[1600] = 4'b1101;
	mem[1601] = 4'b1110;
	mem[1602] = 4'b1111;
	mem[1603] = 4'b1111;
	mem[1604] = 4'b1111;
	mem[1605] = 4'b1110;
	mem[1606] = 4'b1110;
	mem[1607] = 4'b0101;
	mem[1608] = 4'b0001;
	mem[1609] = 4'b0000;
	mem[1610] = 4'b0000;
	mem[1611] = 4'b0000;
	mem[1612] = 4'b0000;
	mem[1613] = 4'b0000;
	mem[1614] = 4'b0000;
	mem[1615] = 4'b0000;
	mem[1616] = 4'b0000;
	mem[1617] = 4'b0000;
	mem[1618] = 4'b0000;
	mem[1619] = 4'b0000;
	mem[1620] = 4'b0000;
	mem[1621] = 4'b0000;
	mem[1622] = 4'b0000;
	mem[1623] = 4'b0000;
	mem[1624] = 4'b0000;
	mem[1625] = 4'b0000;
	mem[1626] = 4'b0000;
	mem[1627] = 4'b0000;
	mem[1628] = 4'b0000;
	mem[1629] = 4'b0000;
	mem[1630] = 4'b0000;
	mem[1631] = 4'b0000;
	mem[1632] = 4'b0000;
	mem[1633] = 4'b0000;
	mem[1634] = 4'b0000;
	mem[1635] = 4'b0000;
	mem[1636] = 4'b0000;
	mem[1637] = 4'b0000;
	mem[1638] = 4'b0000;
	mem[1639] = 4'b0000;
	mem[1640] = 4'b0000;
	mem[1641] = 4'b0000;
	mem[1642] = 4'b0000;
	mem[1643] = 4'b0000;
	mem[1644] = 4'b0000;
	mem[1645] = 4'b0000;
	mem[1646] = 4'b0000;
	mem[1647] = 4'b0000;
	mem[1648] = 4'b0000;
	mem[1649] = 4'b0000;
	mem[1650] = 4'b0000;
	mem[1651] = 4'b0000;
	mem[1652] = 4'b0000;
	mem[1653] = 4'b0000;
	mem[1654] = 4'b0000;
	mem[1655] = 4'b0000;
	mem[1656] = 4'b0000;
	mem[1657] = 4'b0000;
	mem[1658] = 4'b0000;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0111;
	mem[1668] = 4'b1100;
	mem[1669] = 4'b1101;
	mem[1670] = 4'b1101;
	mem[1671] = 4'b1101;
	mem[1672] = 4'b1101;
	mem[1673] = 4'b1101;
	mem[1674] = 4'b1101;
	mem[1675] = 4'b1101;
	mem[1676] = 4'b1101;
	mem[1677] = 4'b1101;
	mem[1678] = 4'b1101;
	mem[1679] = 4'b1101;
	mem[1680] = 4'b1101;
	mem[1681] = 4'b1101;
	mem[1682] = 4'b1101;
	mem[1683] = 4'b1101;
	mem[1684] = 4'b1111;
	mem[1685] = 4'b1111;
	mem[1686] = 4'b1111;
	mem[1687] = 4'b1111;
	mem[1688] = 4'b1111;
	mem[1689] = 4'b1111;
	mem[1690] = 4'b1111;
	mem[1691] = 4'b1111;
	mem[1692] = 4'b1111;
	mem[1693] = 4'b1111;
	mem[1694] = 4'b1111;
	mem[1695] = 4'b1111;
	mem[1696] = 4'b1111;
	mem[1697] = 4'b1111;
	mem[1698] = 4'b1111;
	mem[1699] = 4'b1111;
	mem[1700] = 4'b1111;
	mem[1701] = 4'b1111;
	mem[1702] = 4'b1111;
	mem[1703] = 4'b1111;
	mem[1704] = 4'b1111;
	mem[1705] = 4'b1111;
	mem[1706] = 4'b1111;
	mem[1707] = 4'b1111;
	mem[1708] = 4'b1111;
	mem[1709] = 4'b1111;
	mem[1710] = 4'b1111;
	mem[1711] = 4'b1111;
	mem[1712] = 4'b1111;
	mem[1713] = 4'b1111;
	mem[1714] = 4'b1111;
	mem[1715] = 4'b1111;
	mem[1716] = 4'b1111;
	mem[1717] = 4'b1111;
	mem[1718] = 4'b1111;
	mem[1719] = 4'b1111;
	mem[1720] = 4'b1111;
	mem[1721] = 4'b1111;
	mem[1722] = 4'b1111;
	mem[1723] = 4'b1110;
	mem[1724] = 4'b1111;
	mem[1725] = 4'b1111;
	mem[1726] = 4'b1111;
	mem[1727] = 4'b1111;
	mem[1728] = 4'b1101;
	mem[1729] = 4'b1101;
	mem[1730] = 4'b1110;
	mem[1731] = 4'b1110;
	mem[1732] = 4'b1110;
	mem[1733] = 4'b1101;
	mem[1734] = 4'b1111;
	mem[1735] = 4'b1000;
	mem[1736] = 4'b0101;
	mem[1737] = 4'b0101;
	mem[1738] = 4'b0101;
	mem[1739] = 4'b0101;
	mem[1740] = 4'b0101;
	mem[1741] = 4'b0101;
	mem[1742] = 4'b0101;
	mem[1743] = 4'b0101;
	mem[1744] = 4'b0101;
	mem[1745] = 4'b0101;
	mem[1746] = 4'b0101;
	mem[1747] = 4'b0101;
	mem[1748] = 4'b0101;
	mem[1749] = 4'b0101;
	mem[1750] = 4'b0101;
	mem[1751] = 4'b0101;
	mem[1752] = 4'b0101;
	mem[1753] = 4'b0101;
	mem[1754] = 4'b0101;
	mem[1755] = 4'b0101;
	mem[1756] = 4'b0101;
	mem[1757] = 4'b0101;
	mem[1758] = 4'b0101;
	mem[1759] = 4'b0101;
	mem[1760] = 4'b0101;
	mem[1761] = 4'b0101;
	mem[1762] = 4'b0101;
	mem[1763] = 4'b0101;
	mem[1764] = 4'b0101;
	mem[1765] = 4'b0101;
	mem[1766] = 4'b0101;
	mem[1767] = 4'b0101;
	mem[1768] = 4'b0101;
	mem[1769] = 4'b0101;
	mem[1770] = 4'b0101;
	mem[1771] = 4'b0101;
	mem[1772] = 4'b0101;
	mem[1773] = 4'b0110;
	mem[1774] = 4'b0110;
	mem[1775] = 4'b0110;
	mem[1776] = 4'b0110;
	mem[1777] = 4'b0110;
	mem[1778] = 4'b0101;
	mem[1779] = 4'b0101;
	mem[1780] = 4'b0101;
	mem[1781] = 4'b0101;
	mem[1782] = 4'b0101;
	mem[1783] = 4'b0110;
	mem[1784] = 4'b0000;
	mem[1785] = 4'b0000;
	mem[1786] = 4'b0000;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0111;
	mem[1796] = 4'b1100;
	mem[1797] = 4'b1101;
	mem[1798] = 4'b1101;
	mem[1799] = 4'b1101;
	mem[1800] = 4'b1101;
	mem[1801] = 4'b1101;
	mem[1802] = 4'b1101;
	mem[1803] = 4'b1101;
	mem[1804] = 4'b1101;
	mem[1805] = 4'b1101;
	mem[1806] = 4'b1101;
	mem[1807] = 4'b1101;
	mem[1808] = 4'b1101;
	mem[1809] = 4'b1101;
	mem[1810] = 4'b1101;
	mem[1811] = 4'b1101;
	mem[1812] = 4'b1111;
	mem[1813] = 4'b1111;
	mem[1814] = 4'b1111;
	mem[1815] = 4'b1111;
	mem[1816] = 4'b1111;
	mem[1817] = 4'b1111;
	mem[1818] = 4'b1111;
	mem[1819] = 4'b1111;
	mem[1820] = 4'b1111;
	mem[1821] = 4'b1111;
	mem[1822] = 4'b1111;
	mem[1823] = 4'b1111;
	mem[1824] = 4'b1111;
	mem[1825] = 4'b1111;
	mem[1826] = 4'b1111;
	mem[1827] = 4'b1111;
	mem[1828] = 4'b1111;
	mem[1829] = 4'b1111;
	mem[1830] = 4'b1111;
	mem[1831] = 4'b1111;
	mem[1832] = 4'b1111;
	mem[1833] = 4'b1111;
	mem[1834] = 4'b1111;
	mem[1835] = 4'b1111;
	mem[1836] = 4'b1111;
	mem[1837] = 4'b1111;
	mem[1838] = 4'b1111;
	mem[1839] = 4'b1111;
	mem[1840] = 4'b1111;
	mem[1841] = 4'b1111;
	mem[1842] = 4'b1111;
	mem[1843] = 4'b1111;
	mem[1844] = 4'b1111;
	mem[1845] = 4'b1111;
	mem[1846] = 4'b1111;
	mem[1847] = 4'b1111;
	mem[1848] = 4'b1111;
	mem[1849] = 4'b1110;
	mem[1850] = 4'b1101;
	mem[1851] = 4'b1101;
	mem[1852] = 4'b1101;
	mem[1853] = 4'b1110;
	mem[1854] = 4'b1111;
	mem[1855] = 4'b1111;
	mem[1856] = 4'b1111;
	mem[1857] = 4'b1101;
	mem[1858] = 4'b1101;
	mem[1859] = 4'b1101;
	mem[1860] = 4'b1101;
	mem[1861] = 4'b1110;
	mem[1862] = 4'b1111;
	mem[1863] = 4'b1000;
	mem[1864] = 4'b0101;
	mem[1865] = 4'b0110;
	mem[1866] = 4'b0110;
	mem[1867] = 4'b0110;
	mem[1868] = 4'b0110;
	mem[1869] = 4'b0110;
	mem[1870] = 4'b0110;
	mem[1871] = 4'b0110;
	mem[1872] = 4'b0110;
	mem[1873] = 4'b0110;
	mem[1874] = 4'b0110;
	mem[1875] = 4'b0110;
	mem[1876] = 4'b0110;
	mem[1877] = 4'b0110;
	mem[1878] = 4'b0110;
	mem[1879] = 4'b0110;
	mem[1880] = 4'b0110;
	mem[1881] = 4'b0110;
	mem[1882] = 4'b0110;
	mem[1883] = 4'b0110;
	mem[1884] = 4'b0110;
	mem[1885] = 4'b0110;
	mem[1886] = 4'b0110;
	mem[1887] = 4'b0110;
	mem[1888] = 4'b0110;
	mem[1889] = 4'b0110;
	mem[1890] = 4'b0110;
	mem[1891] = 4'b0110;
	mem[1892] = 4'b0110;
	mem[1893] = 4'b0110;
	mem[1894] = 4'b0110;
	mem[1895] = 4'b0110;
	mem[1896] = 4'b0110;
	mem[1897] = 4'b0110;
	mem[1898] = 4'b0110;
	mem[1899] = 4'b0110;
	mem[1900] = 4'b0110;
	mem[1901] = 4'b0111;
	mem[1902] = 4'b0111;
	mem[1903] = 4'b0110;
	mem[1904] = 4'b0110;
	mem[1905] = 4'b0111;
	mem[1906] = 4'b0111;
	mem[1907] = 4'b0110;
	mem[1908] = 4'b0110;
	mem[1909] = 4'b0110;
	mem[1910] = 4'b0110;
	mem[1911] = 4'b0110;
	mem[1912] = 4'b0000;
	mem[1913] = 4'b0000;
	mem[1914] = 4'b0000;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0111;
	mem[1924] = 4'b1100;
	mem[1925] = 4'b1101;
	mem[1926] = 4'b1101;
	mem[1927] = 4'b1101;
	mem[1928] = 4'b1101;
	mem[1929] = 4'b1101;
	mem[1930] = 4'b1101;
	mem[1931] = 4'b1101;
	mem[1932] = 4'b1101;
	mem[1933] = 4'b1101;
	mem[1934] = 4'b1101;
	mem[1935] = 4'b1101;
	mem[1936] = 4'b1101;
	mem[1937] = 4'b1101;
	mem[1938] = 4'b1101;
	mem[1939] = 4'b1101;
	mem[1940] = 4'b1111;
	mem[1941] = 4'b1111;
	mem[1942] = 4'b1111;
	mem[1943] = 4'b1111;
	mem[1944] = 4'b1111;
	mem[1945] = 4'b1111;
	mem[1946] = 4'b1111;
	mem[1947] = 4'b1111;
	mem[1948] = 4'b1111;
	mem[1949] = 4'b1111;
	mem[1950] = 4'b1111;
	mem[1951] = 4'b1111;
	mem[1952] = 4'b1111;
	mem[1953] = 4'b1111;
	mem[1954] = 4'b1111;
	mem[1955] = 4'b1111;
	mem[1956] = 4'b1111;
	mem[1957] = 4'b1111;
	mem[1958] = 4'b1111;
	mem[1959] = 4'b1111;
	mem[1960] = 4'b1111;
	mem[1961] = 4'b1111;
	mem[1962] = 4'b1111;
	mem[1963] = 4'b1111;
	mem[1964] = 4'b1111;
	mem[1965] = 4'b1111;
	mem[1966] = 4'b1111;
	mem[1967] = 4'b1111;
	mem[1968] = 4'b1111;
	mem[1969] = 4'b1111;
	mem[1970] = 4'b1111;
	mem[1971] = 4'b1111;
	mem[1972] = 4'b1111;
	mem[1973] = 4'b1111;
	mem[1974] = 4'b1111;
	mem[1975] = 4'b1111;
	mem[1976] = 4'b1111;
	mem[1977] = 4'b1101;
	mem[1978] = 4'b1110;
	mem[1979] = 4'b1110;
	mem[1980] = 4'b1101;
	mem[1981] = 4'b1101;
	mem[1982] = 4'b1110;
	mem[1983] = 4'b1111;
	mem[1984] = 4'b1111;
	mem[1985] = 4'b1111;
	mem[1986] = 4'b1111;
	mem[1987] = 4'b1111;
	mem[1988] = 4'b1111;
	mem[1989] = 4'b1111;
	mem[1990] = 4'b1111;
	mem[1991] = 4'b1000;
	mem[1992] = 4'b0110;
	mem[1993] = 4'b0110;
	mem[1994] = 4'b0110;
	mem[1995] = 4'b0110;
	mem[1996] = 4'b0110;
	mem[1997] = 4'b0110;
	mem[1998] = 4'b0110;
	mem[1999] = 4'b0110;
	mem[2000] = 4'b0110;
	mem[2001] = 4'b0110;
	mem[2002] = 4'b0110;
	mem[2003] = 4'b0110;
	mem[2004] = 4'b0110;
	mem[2005] = 4'b0110;
	mem[2006] = 4'b0110;
	mem[2007] = 4'b0110;
	mem[2008] = 4'b0110;
	mem[2009] = 4'b0110;
	mem[2010] = 4'b0110;
	mem[2011] = 4'b0110;
	mem[2012] = 4'b0110;
	mem[2013] = 4'b0110;
	mem[2014] = 4'b0110;
	mem[2015] = 4'b0110;
	mem[2016] = 4'b0110;
	mem[2017] = 4'b0110;
	mem[2018] = 4'b0110;
	mem[2019] = 4'b0110;
	mem[2020] = 4'b0110;
	mem[2021] = 4'b0110;
	mem[2022] = 4'b0110;
	mem[2023] = 4'b0110;
	mem[2024] = 4'b0110;
	mem[2025] = 4'b0110;
	mem[2026] = 4'b0110;
	mem[2027] = 4'b0110;
	mem[2028] = 4'b0111;
	mem[2029] = 4'b0111;
	mem[2030] = 4'b0110;
	mem[2031] = 4'b0110;
	mem[2032] = 4'b0110;
	mem[2033] = 4'b0110;
	mem[2034] = 4'b0110;
	mem[2035] = 4'b0111;
	mem[2036] = 4'b0110;
	mem[2037] = 4'b0110;
	mem[2038] = 4'b0110;
	mem[2039] = 4'b0110;
	mem[2040] = 4'b0000;
	mem[2041] = 4'b0000;
	mem[2042] = 4'b0000;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0111;
	mem[2052] = 4'b1100;
	mem[2053] = 4'b1101;
	mem[2054] = 4'b1101;
	mem[2055] = 4'b1101;
	mem[2056] = 4'b1101;
	mem[2057] = 4'b1101;
	mem[2058] = 4'b1101;
	mem[2059] = 4'b1101;
	mem[2060] = 4'b1101;
	mem[2061] = 4'b1101;
	mem[2062] = 4'b1101;
	mem[2063] = 4'b1101;
	mem[2064] = 4'b1101;
	mem[2065] = 4'b1101;
	mem[2066] = 4'b1101;
	mem[2067] = 4'b1101;
	mem[2068] = 4'b1111;
	mem[2069] = 4'b1111;
	mem[2070] = 4'b1111;
	mem[2071] = 4'b1111;
	mem[2072] = 4'b1111;
	mem[2073] = 4'b1111;
	mem[2074] = 4'b1111;
	mem[2075] = 4'b1111;
	mem[2076] = 4'b1111;
	mem[2077] = 4'b1111;
	mem[2078] = 4'b1111;
	mem[2079] = 4'b1111;
	mem[2080] = 4'b1111;
	mem[2081] = 4'b1111;
	mem[2082] = 4'b1111;
	mem[2083] = 4'b1111;
	mem[2084] = 4'b1111;
	mem[2085] = 4'b1111;
	mem[2086] = 4'b1111;
	mem[2087] = 4'b1111;
	mem[2088] = 4'b1111;
	mem[2089] = 4'b1111;
	mem[2090] = 4'b1111;
	mem[2091] = 4'b1111;
	mem[2092] = 4'b1111;
	mem[2093] = 4'b1111;
	mem[2094] = 4'b1111;
	mem[2095] = 4'b1111;
	mem[2096] = 4'b1111;
	mem[2097] = 4'b1111;
	mem[2098] = 4'b1111;
	mem[2099] = 4'b1111;
	mem[2100] = 4'b1111;
	mem[2101] = 4'b1111;
	mem[2102] = 4'b1111;
	mem[2103] = 4'b1111;
	mem[2104] = 4'b1110;
	mem[2105] = 4'b1110;
	mem[2106] = 4'b1111;
	mem[2107] = 4'b1111;
	mem[2108] = 4'b1111;
	mem[2109] = 4'b1101;
	mem[2110] = 4'b1101;
	mem[2111] = 4'b1110;
	mem[2112] = 4'b1111;
	mem[2113] = 4'b1111;
	mem[2114] = 4'b1111;
	mem[2115] = 4'b1111;
	mem[2116] = 4'b1111;
	mem[2117] = 4'b1111;
	mem[2118] = 4'b1111;
	mem[2119] = 4'b1000;
	mem[2120] = 4'b0110;
	mem[2121] = 4'b0110;
	mem[2122] = 4'b0110;
	mem[2123] = 4'b0110;
	mem[2124] = 4'b0110;
	mem[2125] = 4'b0110;
	mem[2126] = 4'b0110;
	mem[2127] = 4'b0110;
	mem[2128] = 4'b0110;
	mem[2129] = 4'b0110;
	mem[2130] = 4'b0110;
	mem[2131] = 4'b0110;
	mem[2132] = 4'b0110;
	mem[2133] = 4'b0110;
	mem[2134] = 4'b0110;
	mem[2135] = 4'b0110;
	mem[2136] = 4'b0110;
	mem[2137] = 4'b0110;
	mem[2138] = 4'b0110;
	mem[2139] = 4'b0110;
	mem[2140] = 4'b0110;
	mem[2141] = 4'b0110;
	mem[2142] = 4'b0110;
	mem[2143] = 4'b0110;
	mem[2144] = 4'b0110;
	mem[2145] = 4'b0110;
	mem[2146] = 4'b0110;
	mem[2147] = 4'b0110;
	mem[2148] = 4'b0110;
	mem[2149] = 4'b0110;
	mem[2150] = 4'b0110;
	mem[2151] = 4'b0110;
	mem[2152] = 4'b0110;
	mem[2153] = 4'b0110;
	mem[2154] = 4'b0110;
	mem[2155] = 4'b0110;
	mem[2156] = 4'b0111;
	mem[2157] = 4'b0111;
	mem[2158] = 4'b0110;
	mem[2159] = 4'b0110;
	mem[2160] = 4'b0110;
	mem[2161] = 4'b0111;
	mem[2162] = 4'b0111;
	mem[2163] = 4'b0111;
	mem[2164] = 4'b0111;
	mem[2165] = 4'b0110;
	mem[2166] = 4'b0110;
	mem[2167] = 4'b0110;
	mem[2168] = 4'b0000;
	mem[2169] = 4'b0000;
	mem[2170] = 4'b0000;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0111;
	mem[2180] = 4'b1100;
	mem[2181] = 4'b1101;
	mem[2182] = 4'b1101;
	mem[2183] = 4'b1101;
	mem[2184] = 4'b1101;
	mem[2185] = 4'b1101;
	mem[2186] = 4'b1101;
	mem[2187] = 4'b1101;
	mem[2188] = 4'b1101;
	mem[2189] = 4'b1101;
	mem[2190] = 4'b1101;
	mem[2191] = 4'b1101;
	mem[2192] = 4'b1101;
	mem[2193] = 4'b1101;
	mem[2194] = 4'b1101;
	mem[2195] = 4'b1101;
	mem[2196] = 4'b1111;
	mem[2197] = 4'b1111;
	mem[2198] = 4'b1111;
	mem[2199] = 4'b1111;
	mem[2200] = 4'b1111;
	mem[2201] = 4'b1111;
	mem[2202] = 4'b1111;
	mem[2203] = 4'b1111;
	mem[2204] = 4'b1111;
	mem[2205] = 4'b1111;
	mem[2206] = 4'b1111;
	mem[2207] = 4'b1111;
	mem[2208] = 4'b1111;
	mem[2209] = 4'b1111;
	mem[2210] = 4'b1111;
	mem[2211] = 4'b1111;
	mem[2212] = 4'b1111;
	mem[2213] = 4'b1111;
	mem[2214] = 4'b1111;
	mem[2215] = 4'b1111;
	mem[2216] = 4'b1111;
	mem[2217] = 4'b1111;
	mem[2218] = 4'b1111;
	mem[2219] = 4'b1111;
	mem[2220] = 4'b1111;
	mem[2221] = 4'b1111;
	mem[2222] = 4'b1111;
	mem[2223] = 4'b1111;
	mem[2224] = 4'b1111;
	mem[2225] = 4'b1111;
	mem[2226] = 4'b1111;
	mem[2227] = 4'b1111;
	mem[2228] = 4'b1111;
	mem[2229] = 4'b1111;
	mem[2230] = 4'b1110;
	mem[2231] = 4'b1101;
	mem[2232] = 4'b1101;
	mem[2233] = 4'b1111;
	mem[2234] = 4'b1111;
	mem[2235] = 4'b1111;
	mem[2236] = 4'b1111;
	mem[2237] = 4'b1111;
	mem[2238] = 4'b1101;
	mem[2239] = 4'b1101;
	mem[2240] = 4'b1110;
	mem[2241] = 4'b1111;
	mem[2242] = 4'b1111;
	mem[2243] = 4'b1111;
	mem[2244] = 4'b1111;
	mem[2245] = 4'b1111;
	mem[2246] = 4'b1111;
	mem[2247] = 4'b1000;
	mem[2248] = 4'b0110;
	mem[2249] = 4'b0110;
	mem[2250] = 4'b0110;
	mem[2251] = 4'b0110;
	mem[2252] = 4'b0110;
	mem[2253] = 4'b0110;
	mem[2254] = 4'b0110;
	mem[2255] = 4'b0110;
	mem[2256] = 4'b0110;
	mem[2257] = 4'b0110;
	mem[2258] = 4'b0110;
	mem[2259] = 4'b0110;
	mem[2260] = 4'b0110;
	mem[2261] = 4'b0110;
	mem[2262] = 4'b0110;
	mem[2263] = 4'b0110;
	mem[2264] = 4'b0110;
	mem[2265] = 4'b0110;
	mem[2266] = 4'b0110;
	mem[2267] = 4'b0110;
	mem[2268] = 4'b0110;
	mem[2269] = 4'b0110;
	mem[2270] = 4'b0110;
	mem[2271] = 4'b0110;
	mem[2272] = 4'b0110;
	mem[2273] = 4'b0110;
	mem[2274] = 4'b0110;
	mem[2275] = 4'b0110;
	mem[2276] = 4'b0110;
	mem[2277] = 4'b0110;
	mem[2278] = 4'b0110;
	mem[2279] = 4'b0110;
	mem[2280] = 4'b0110;
	mem[2281] = 4'b0110;
	mem[2282] = 4'b0110;
	mem[2283] = 4'b0110;
	mem[2284] = 4'b0110;
	mem[2285] = 4'b0111;
	mem[2286] = 4'b0110;
	mem[2287] = 4'b0111;
	mem[2288] = 4'b0111;
	mem[2289] = 4'b0111;
	mem[2290] = 4'b0111;
	mem[2291] = 4'b0111;
	mem[2292] = 4'b0111;
	mem[2293] = 4'b0110;
	mem[2294] = 4'b0110;
	mem[2295] = 4'b0110;
	mem[2296] = 4'b0000;
	mem[2297] = 4'b0000;
	mem[2298] = 4'b0000;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0111;
	mem[2308] = 4'b1100;
	mem[2309] = 4'b1101;
	mem[2310] = 4'b1101;
	mem[2311] = 4'b1101;
	mem[2312] = 4'b1101;
	mem[2313] = 4'b1101;
	mem[2314] = 4'b1101;
	mem[2315] = 4'b1101;
	mem[2316] = 4'b1101;
	mem[2317] = 4'b1101;
	mem[2318] = 4'b1101;
	mem[2319] = 4'b1101;
	mem[2320] = 4'b1101;
	mem[2321] = 4'b1101;
	mem[2322] = 4'b1101;
	mem[2323] = 4'b1101;
	mem[2324] = 4'b1111;
	mem[2325] = 4'b1111;
	mem[2326] = 4'b1111;
	mem[2327] = 4'b1111;
	mem[2328] = 4'b1111;
	mem[2329] = 4'b1111;
	mem[2330] = 4'b1111;
	mem[2331] = 4'b1111;
	mem[2332] = 4'b1111;
	mem[2333] = 4'b1111;
	mem[2334] = 4'b1111;
	mem[2335] = 4'b1111;
	mem[2336] = 4'b1111;
	mem[2337] = 4'b1111;
	mem[2338] = 4'b1111;
	mem[2339] = 4'b1111;
	mem[2340] = 4'b1111;
	mem[2341] = 4'b1111;
	mem[2342] = 4'b1111;
	mem[2343] = 4'b1111;
	mem[2344] = 4'b1111;
	mem[2345] = 4'b1111;
	mem[2346] = 4'b1111;
	mem[2347] = 4'b1111;
	mem[2348] = 4'b1111;
	mem[2349] = 4'b1111;
	mem[2350] = 4'b1111;
	mem[2351] = 4'b1111;
	mem[2352] = 4'b1111;
	mem[2353] = 4'b1111;
	mem[2354] = 4'b1111;
	mem[2355] = 4'b1111;
	mem[2356] = 4'b1111;
	mem[2357] = 4'b1111;
	mem[2358] = 4'b1111;
	mem[2359] = 4'b1101;
	mem[2360] = 4'b1101;
	mem[2361] = 4'b1110;
	mem[2362] = 4'b1111;
	mem[2363] = 4'b1111;
	mem[2364] = 4'b1111;
	mem[2365] = 4'b1111;
	mem[2366] = 4'b1111;
	mem[2367] = 4'b1101;
	mem[2368] = 4'b1101;
	mem[2369] = 4'b1111;
	mem[2370] = 4'b1111;
	mem[2371] = 4'b1111;
	mem[2372] = 4'b1111;
	mem[2373] = 4'b1111;
	mem[2374] = 4'b1111;
	mem[2375] = 4'b1000;
	mem[2376] = 4'b0110;
	mem[2377] = 4'b0110;
	mem[2378] = 4'b0110;
	mem[2379] = 4'b0110;
	mem[2380] = 4'b0110;
	mem[2381] = 4'b0110;
	mem[2382] = 4'b0110;
	mem[2383] = 4'b0110;
	mem[2384] = 4'b0110;
	mem[2385] = 4'b0110;
	mem[2386] = 4'b0110;
	mem[2387] = 4'b0110;
	mem[2388] = 4'b0110;
	mem[2389] = 4'b0110;
	mem[2390] = 4'b0110;
	mem[2391] = 4'b0110;
	mem[2392] = 4'b0110;
	mem[2393] = 4'b0110;
	mem[2394] = 4'b0110;
	mem[2395] = 4'b0110;
	mem[2396] = 4'b0110;
	mem[2397] = 4'b0110;
	mem[2398] = 4'b0110;
	mem[2399] = 4'b0110;
	mem[2400] = 4'b0110;
	mem[2401] = 4'b0110;
	mem[2402] = 4'b0110;
	mem[2403] = 4'b0110;
	mem[2404] = 4'b0110;
	mem[2405] = 4'b0110;
	mem[2406] = 4'b0110;
	mem[2407] = 4'b0110;
	mem[2408] = 4'b0110;
	mem[2409] = 4'b0110;
	mem[2410] = 4'b0110;
	mem[2411] = 4'b0110;
	mem[2412] = 4'b0110;
	mem[2413] = 4'b0111;
	mem[2414] = 4'b0111;
	mem[2415] = 4'b0111;
	mem[2416] = 4'b0111;
	mem[2417] = 4'b0111;
	mem[2418] = 4'b0111;
	mem[2419] = 4'b0111;
	mem[2420] = 4'b0111;
	mem[2421] = 4'b0110;
	mem[2422] = 4'b0110;
	mem[2423] = 4'b0110;
	mem[2424] = 4'b0000;
	mem[2425] = 4'b0000;
	mem[2426] = 4'b0001;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0111;
	mem[2436] = 4'b1100;
	mem[2437] = 4'b1101;
	mem[2438] = 4'b1101;
	mem[2439] = 4'b1101;
	mem[2440] = 4'b1101;
	mem[2441] = 4'b1101;
	mem[2442] = 4'b1101;
	mem[2443] = 4'b1101;
	mem[2444] = 4'b1101;
	mem[2445] = 4'b1101;
	mem[2446] = 4'b1101;
	mem[2447] = 4'b1101;
	mem[2448] = 4'b1101;
	mem[2449] = 4'b1101;
	mem[2450] = 4'b1101;
	mem[2451] = 4'b1101;
	mem[2452] = 4'b1111;
	mem[2453] = 4'b1111;
	mem[2454] = 4'b1111;
	mem[2455] = 4'b1111;
	mem[2456] = 4'b1111;
	mem[2457] = 4'b1111;
	mem[2458] = 4'b1111;
	mem[2459] = 4'b1111;
	mem[2460] = 4'b1111;
	mem[2461] = 4'b1111;
	mem[2462] = 4'b1111;
	mem[2463] = 4'b1111;
	mem[2464] = 4'b1111;
	mem[2465] = 4'b1111;
	mem[2466] = 4'b1111;
	mem[2467] = 4'b1111;
	mem[2468] = 4'b1111;
	mem[2469] = 4'b1111;
	mem[2470] = 4'b1111;
	mem[2471] = 4'b1111;
	mem[2472] = 4'b1111;
	mem[2473] = 4'b1111;
	mem[2474] = 4'b1111;
	mem[2475] = 4'b1111;
	mem[2476] = 4'b1111;
	mem[2477] = 4'b1111;
	mem[2478] = 4'b1111;
	mem[2479] = 4'b1111;
	mem[2480] = 4'b1111;
	mem[2481] = 4'b1111;
	mem[2482] = 4'b1111;
	mem[2483] = 4'b1111;
	mem[2484] = 4'b1111;
	mem[2485] = 4'b1111;
	mem[2486] = 4'b1111;
	mem[2487] = 4'b1111;
	mem[2488] = 4'b1101;
	mem[2489] = 4'b1101;
	mem[2490] = 4'b1110;
	mem[2491] = 4'b1111;
	mem[2492] = 4'b1111;
	mem[2493] = 4'b1111;
	mem[2494] = 4'b1111;
	mem[2495] = 4'b1111;
	mem[2496] = 4'b1110;
	mem[2497] = 4'b1111;
	mem[2498] = 4'b1111;
	mem[2499] = 4'b1111;
	mem[2500] = 4'b1111;
	mem[2501] = 4'b1111;
	mem[2502] = 4'b1111;
	mem[2503] = 4'b1000;
	mem[2504] = 4'b0110;
	mem[2505] = 4'b0110;
	mem[2506] = 4'b0110;
	mem[2507] = 4'b0110;
	mem[2508] = 4'b0110;
	mem[2509] = 4'b0110;
	mem[2510] = 4'b0110;
	mem[2511] = 4'b0110;
	mem[2512] = 4'b0110;
	mem[2513] = 4'b0110;
	mem[2514] = 4'b0110;
	mem[2515] = 4'b0110;
	mem[2516] = 4'b0110;
	mem[2517] = 4'b0110;
	mem[2518] = 4'b0110;
	mem[2519] = 4'b0110;
	mem[2520] = 4'b0110;
	mem[2521] = 4'b0110;
	mem[2522] = 4'b0110;
	mem[2523] = 4'b0110;
	mem[2524] = 4'b0110;
	mem[2525] = 4'b0110;
	mem[2526] = 4'b0110;
	mem[2527] = 4'b0110;
	mem[2528] = 4'b0110;
	mem[2529] = 4'b0110;
	mem[2530] = 4'b0110;
	mem[2531] = 4'b0110;
	mem[2532] = 4'b0110;
	mem[2533] = 4'b0110;
	mem[2534] = 4'b0110;
	mem[2535] = 4'b0110;
	mem[2536] = 4'b0110;
	mem[2537] = 4'b0110;
	mem[2538] = 4'b0110;
	mem[2539] = 4'b0110;
	mem[2540] = 4'b0110;
	mem[2541] = 4'b0110;
	mem[2542] = 4'b0111;
	mem[2543] = 4'b0111;
	mem[2544] = 4'b0111;
	mem[2545] = 4'b0111;
	mem[2546] = 4'b0111;
	mem[2547] = 4'b0111;
	mem[2548] = 4'b0111;
	mem[2549] = 4'b0110;
	mem[2550] = 4'b0110;
	mem[2551] = 4'b0111;
	mem[2552] = 4'b0001;
	mem[2553] = 4'b0001;
	mem[2554] = 4'b0000;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b0111;
	mem[2564] = 4'b1100;
	mem[2565] = 4'b1101;
	mem[2566] = 4'b1101;
	mem[2567] = 4'b1101;
	mem[2568] = 4'b1101;
	mem[2569] = 4'b1101;
	mem[2570] = 4'b1101;
	mem[2571] = 4'b1101;
	mem[2572] = 4'b1101;
	mem[2573] = 4'b1101;
	mem[2574] = 4'b1101;
	mem[2575] = 4'b1101;
	mem[2576] = 4'b1101;
	mem[2577] = 4'b1101;
	mem[2578] = 4'b1101;
	mem[2579] = 4'b1101;
	mem[2580] = 4'b1111;
	mem[2581] = 4'b1111;
	mem[2582] = 4'b1111;
	mem[2583] = 4'b1111;
	mem[2584] = 4'b1111;
	mem[2585] = 4'b1111;
	mem[2586] = 4'b1111;
	mem[2587] = 4'b1111;
	mem[2588] = 4'b1111;
	mem[2589] = 4'b1111;
	mem[2590] = 4'b1111;
	mem[2591] = 4'b1111;
	mem[2592] = 4'b1111;
	mem[2593] = 4'b1111;
	mem[2594] = 4'b1111;
	mem[2595] = 4'b1111;
	mem[2596] = 4'b1111;
	mem[2597] = 4'b1111;
	mem[2598] = 4'b1111;
	mem[2599] = 4'b1111;
	mem[2600] = 4'b1111;
	mem[2601] = 4'b1111;
	mem[2602] = 4'b1111;
	mem[2603] = 4'b1111;
	mem[2604] = 4'b1111;
	mem[2605] = 4'b1111;
	mem[2606] = 4'b1111;
	mem[2607] = 4'b1111;
	mem[2608] = 4'b1111;
	mem[2609] = 4'b1111;
	mem[2610] = 4'b1111;
	mem[2611] = 4'b1111;
	mem[2612] = 4'b1110;
	mem[2613] = 4'b1111;
	mem[2614] = 4'b1111;
	mem[2615] = 4'b1111;
	mem[2616] = 4'b1111;
	mem[2617] = 4'b1101;
	mem[2618] = 4'b1101;
	mem[2619] = 4'b1110;
	mem[2620] = 4'b1111;
	mem[2621] = 4'b1111;
	mem[2622] = 4'b1111;
	mem[2623] = 4'b1111;
	mem[2624] = 4'b1111;
	mem[2625] = 4'b1111;
	mem[2626] = 4'b1111;
	mem[2627] = 4'b1111;
	mem[2628] = 4'b1111;
	mem[2629] = 4'b1111;
	mem[2630] = 4'b1111;
	mem[2631] = 4'b1000;
	mem[2632] = 4'b0110;
	mem[2633] = 4'b0110;
	mem[2634] = 4'b0110;
	mem[2635] = 4'b0110;
	mem[2636] = 4'b0110;
	mem[2637] = 4'b0110;
	mem[2638] = 4'b0110;
	mem[2639] = 4'b0110;
	mem[2640] = 4'b0110;
	mem[2641] = 4'b0110;
	mem[2642] = 4'b0110;
	mem[2643] = 4'b0110;
	mem[2644] = 4'b0110;
	mem[2645] = 4'b0110;
	mem[2646] = 4'b0110;
	mem[2647] = 4'b0110;
	mem[2648] = 4'b0110;
	mem[2649] = 4'b0110;
	mem[2650] = 4'b0110;
	mem[2651] = 4'b0110;
	mem[2652] = 4'b0110;
	mem[2653] = 4'b0110;
	mem[2654] = 4'b0110;
	mem[2655] = 4'b0110;
	mem[2656] = 4'b0110;
	mem[2657] = 4'b0110;
	mem[2658] = 4'b0110;
	mem[2659] = 4'b0110;
	mem[2660] = 4'b0110;
	mem[2661] = 4'b0110;
	mem[2662] = 4'b0110;
	mem[2663] = 4'b0110;
	mem[2664] = 4'b0110;
	mem[2665] = 4'b0111;
	mem[2666] = 4'b0110;
	mem[2667] = 4'b0110;
	mem[2668] = 4'b0110;
	mem[2669] = 4'b0110;
	mem[2670] = 4'b0110;
	mem[2671] = 4'b0111;
	mem[2672] = 4'b0111;
	mem[2673] = 4'b0111;
	mem[2674] = 4'b0111;
	mem[2675] = 4'b0111;
	mem[2676] = 4'b0110;
	mem[2677] = 4'b0110;
	mem[2678] = 4'b0110;
	mem[2679] = 4'b1000;
	mem[2680] = 4'b0000;
	mem[2681] = 4'b0000;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b0111;
	mem[2692] = 4'b1100;
	mem[2693] = 4'b1101;
	mem[2694] = 4'b1101;
	mem[2695] = 4'b1101;
	mem[2696] = 4'b1101;
	mem[2697] = 4'b1101;
	mem[2698] = 4'b1101;
	mem[2699] = 4'b1101;
	mem[2700] = 4'b1101;
	mem[2701] = 4'b1101;
	mem[2702] = 4'b1101;
	mem[2703] = 4'b1101;
	mem[2704] = 4'b1101;
	mem[2705] = 4'b1101;
	mem[2706] = 4'b1101;
	mem[2707] = 4'b1101;
	mem[2708] = 4'b1111;
	mem[2709] = 4'b1111;
	mem[2710] = 4'b1111;
	mem[2711] = 4'b1111;
	mem[2712] = 4'b1111;
	mem[2713] = 4'b1111;
	mem[2714] = 4'b1111;
	mem[2715] = 4'b1111;
	mem[2716] = 4'b1111;
	mem[2717] = 4'b1111;
	mem[2718] = 4'b1111;
	mem[2719] = 4'b1111;
	mem[2720] = 4'b1111;
	mem[2721] = 4'b1111;
	mem[2722] = 4'b1111;
	mem[2723] = 4'b1111;
	mem[2724] = 4'b1111;
	mem[2725] = 4'b1111;
	mem[2726] = 4'b1111;
	mem[2727] = 4'b1111;
	mem[2728] = 4'b1111;
	mem[2729] = 4'b1111;
	mem[2730] = 4'b1111;
	mem[2731] = 4'b1111;
	mem[2732] = 4'b1111;
	mem[2733] = 4'b1111;
	mem[2734] = 4'b1111;
	mem[2735] = 4'b1111;
	mem[2736] = 4'b1111;
	mem[2737] = 4'b1111;
	mem[2738] = 4'b1110;
	mem[2739] = 4'b1101;
	mem[2740] = 4'b1101;
	mem[2741] = 4'b1101;
	mem[2742] = 4'b1111;
	mem[2743] = 4'b1111;
	mem[2744] = 4'b1111;
	mem[2745] = 4'b1111;
	mem[2746] = 4'b1101;
	mem[2747] = 4'b1101;
	mem[2748] = 4'b1110;
	mem[2749] = 4'b1111;
	mem[2750] = 4'b1111;
	mem[2751] = 4'b1111;
	mem[2752] = 4'b1111;
	mem[2753] = 4'b1111;
	mem[2754] = 4'b1111;
	mem[2755] = 4'b1111;
	mem[2756] = 4'b1111;
	mem[2757] = 4'b1111;
	mem[2758] = 4'b1111;
	mem[2759] = 4'b1000;
	mem[2760] = 4'b0110;
	mem[2761] = 4'b0110;
	mem[2762] = 4'b0110;
	mem[2763] = 4'b0110;
	mem[2764] = 4'b0110;
	mem[2765] = 4'b0110;
	mem[2766] = 4'b0110;
	mem[2767] = 4'b0110;
	mem[2768] = 4'b0110;
	mem[2769] = 4'b0110;
	mem[2770] = 4'b0110;
	mem[2771] = 4'b0110;
	mem[2772] = 4'b0110;
	mem[2773] = 4'b0110;
	mem[2774] = 4'b0110;
	mem[2775] = 4'b0110;
	mem[2776] = 4'b0110;
	mem[2777] = 4'b0110;
	mem[2778] = 4'b0110;
	mem[2779] = 4'b0110;
	mem[2780] = 4'b0110;
	mem[2781] = 4'b0110;
	mem[2782] = 4'b0110;
	mem[2783] = 4'b0110;
	mem[2784] = 4'b0110;
	mem[2785] = 4'b0110;
	mem[2786] = 4'b0110;
	mem[2787] = 4'b0110;
	mem[2788] = 4'b0110;
	mem[2789] = 4'b0111;
	mem[2790] = 4'b0111;
	mem[2791] = 4'b0110;
	mem[2792] = 4'b0111;
	mem[2793] = 4'b0111;
	mem[2794] = 4'b0111;
	mem[2795] = 4'b0110;
	mem[2796] = 4'b0110;
	mem[2797] = 4'b0110;
	mem[2798] = 4'b0110;
	mem[2799] = 4'b0110;
	mem[2800] = 4'b0110;
	mem[2801] = 4'b0110;
	mem[2802] = 4'b0110;
	mem[2803] = 4'b0110;
	mem[2804] = 4'b0110;
	mem[2805] = 4'b0110;
	mem[2806] = 4'b0111;
	mem[2807] = 4'b1000;
	mem[2808] = 4'b0000;
	mem[2809] = 4'b0000;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b0111;
	mem[2820] = 4'b1100;
	mem[2821] = 4'b1101;
	mem[2822] = 4'b1101;
	mem[2823] = 4'b1101;
	mem[2824] = 4'b1101;
	mem[2825] = 4'b1101;
	mem[2826] = 4'b1101;
	mem[2827] = 4'b1101;
	mem[2828] = 4'b1101;
	mem[2829] = 4'b1101;
	mem[2830] = 4'b1101;
	mem[2831] = 4'b1101;
	mem[2832] = 4'b1101;
	mem[2833] = 4'b1101;
	mem[2834] = 4'b1101;
	mem[2835] = 4'b1101;
	mem[2836] = 4'b1111;
	mem[2837] = 4'b1111;
	mem[2838] = 4'b1111;
	mem[2839] = 4'b1111;
	mem[2840] = 4'b1111;
	mem[2841] = 4'b1111;
	mem[2842] = 4'b1111;
	mem[2843] = 4'b1111;
	mem[2844] = 4'b1111;
	mem[2845] = 4'b1111;
	mem[2846] = 4'b1111;
	mem[2847] = 4'b1111;
	mem[2848] = 4'b1111;
	mem[2849] = 4'b1111;
	mem[2850] = 4'b1111;
	mem[2851] = 4'b1111;
	mem[2852] = 4'b1111;
	mem[2853] = 4'b1111;
	mem[2854] = 4'b1111;
	mem[2855] = 4'b1111;
	mem[2856] = 4'b1111;
	mem[2857] = 4'b1111;
	mem[2858] = 4'b1111;
	mem[2859] = 4'b1111;
	mem[2860] = 4'b1111;
	mem[2861] = 4'b1111;
	mem[2862] = 4'b1111;
	mem[2863] = 4'b1111;
	mem[2864] = 4'b1111;
	mem[2865] = 4'b1110;
	mem[2866] = 4'b1101;
	mem[2867] = 4'b1110;
	mem[2868] = 4'b1110;
	mem[2869] = 4'b1101;
	mem[2870] = 4'b1101;
	mem[2871] = 4'b1111;
	mem[2872] = 4'b1111;
	mem[2873] = 4'b1111;
	mem[2874] = 4'b1111;
	mem[2875] = 4'b1101;
	mem[2876] = 4'b1101;
	mem[2877] = 4'b1111;
	mem[2878] = 4'b1111;
	mem[2879] = 4'b1111;
	mem[2880] = 4'b1111;
	mem[2881] = 4'b1111;
	mem[2882] = 4'b1111;
	mem[2883] = 4'b1111;
	mem[2884] = 4'b1111;
	mem[2885] = 4'b1111;
	mem[2886] = 4'b1111;
	mem[2887] = 4'b1000;
	mem[2888] = 4'b0110;
	mem[2889] = 4'b0110;
	mem[2890] = 4'b0110;
	mem[2891] = 4'b0110;
	mem[2892] = 4'b0110;
	mem[2893] = 4'b0110;
	mem[2894] = 4'b0110;
	mem[2895] = 4'b0110;
	mem[2896] = 4'b0110;
	mem[2897] = 4'b0110;
	mem[2898] = 4'b0110;
	mem[2899] = 4'b0110;
	mem[2900] = 4'b0110;
	mem[2901] = 4'b0110;
	mem[2902] = 4'b0110;
	mem[2903] = 4'b0110;
	mem[2904] = 4'b0110;
	mem[2905] = 4'b0110;
	mem[2906] = 4'b0110;
	mem[2907] = 4'b0110;
	mem[2908] = 4'b0110;
	mem[2909] = 4'b0110;
	mem[2910] = 4'b0110;
	mem[2911] = 4'b0110;
	mem[2912] = 4'b0110;
	mem[2913] = 4'b0110;
	mem[2914] = 4'b0110;
	mem[2915] = 4'b0110;
	mem[2916] = 4'b0110;
	mem[2917] = 4'b0110;
	mem[2918] = 4'b0111;
	mem[2919] = 4'b0111;
	mem[2920] = 4'b0111;
	mem[2921] = 4'b0111;
	mem[2922] = 4'b0111;
	mem[2923] = 4'b0111;
	mem[2924] = 4'b0110;
	mem[2925] = 4'b0110;
	mem[2926] = 4'b0110;
	mem[2927] = 4'b0110;
	mem[2928] = 4'b0110;
	mem[2929] = 4'b0110;
	mem[2930] = 4'b0110;
	mem[2931] = 4'b0110;
	mem[2932] = 4'b0110;
	mem[2933] = 4'b0110;
	mem[2934] = 4'b1000;
	mem[2935] = 4'b0111;
	mem[2936] = 4'b0000;
	mem[2937] = 4'b0000;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b0111;
	mem[2948] = 4'b1100;
	mem[2949] = 4'b1101;
	mem[2950] = 4'b1101;
	mem[2951] = 4'b1101;
	mem[2952] = 4'b1101;
	mem[2953] = 4'b1101;
	mem[2954] = 4'b1101;
	mem[2955] = 4'b1101;
	mem[2956] = 4'b1101;
	mem[2957] = 4'b1101;
	mem[2958] = 4'b1101;
	mem[2959] = 4'b1101;
	mem[2960] = 4'b1101;
	mem[2961] = 4'b1101;
	mem[2962] = 4'b1101;
	mem[2963] = 4'b1101;
	mem[2964] = 4'b1111;
	mem[2965] = 4'b1111;
	mem[2966] = 4'b1111;
	mem[2967] = 4'b1111;
	mem[2968] = 4'b1111;
	mem[2969] = 4'b1111;
	mem[2970] = 4'b1111;
	mem[2971] = 4'b1111;
	mem[2972] = 4'b1111;
	mem[2973] = 4'b1111;
	mem[2974] = 4'b1111;
	mem[2975] = 4'b1111;
	mem[2976] = 4'b1111;
	mem[2977] = 4'b1111;
	mem[2978] = 4'b1111;
	mem[2979] = 4'b1111;
	mem[2980] = 4'b1111;
	mem[2981] = 4'b1111;
	mem[2982] = 4'b1111;
	mem[2983] = 4'b1111;
	mem[2984] = 4'b1111;
	mem[2985] = 4'b1111;
	mem[2986] = 4'b1111;
	mem[2987] = 4'b1111;
	mem[2988] = 4'b1111;
	mem[2989] = 4'b1111;
	mem[2990] = 4'b1111;
	mem[2991] = 4'b1111;
	mem[2992] = 4'b1111;
	mem[2993] = 4'b1101;
	mem[2994] = 4'b1110;
	mem[2995] = 4'b1111;
	mem[2996] = 4'b1111;
	mem[2997] = 4'b1101;
	mem[2998] = 4'b1101;
	mem[2999] = 4'b1101;
	mem[3000] = 4'b1111;
	mem[3001] = 4'b1111;
	mem[3002] = 4'b1111;
	mem[3003] = 4'b1111;
	mem[3004] = 4'b1110;
	mem[3005] = 4'b1111;
	mem[3006] = 4'b1111;
	mem[3007] = 4'b1111;
	mem[3008] = 4'b1111;
	mem[3009] = 4'b1111;
	mem[3010] = 4'b1111;
	mem[3011] = 4'b1111;
	mem[3012] = 4'b1111;
	mem[3013] = 4'b1111;
	mem[3014] = 4'b1111;
	mem[3015] = 4'b1000;
	mem[3016] = 4'b0110;
	mem[3017] = 4'b0110;
	mem[3018] = 4'b0110;
	mem[3019] = 4'b0110;
	mem[3020] = 4'b0110;
	mem[3021] = 4'b0110;
	mem[3022] = 4'b0110;
	mem[3023] = 4'b0110;
	mem[3024] = 4'b0110;
	mem[3025] = 4'b0110;
	mem[3026] = 4'b0110;
	mem[3027] = 4'b0110;
	mem[3028] = 4'b0110;
	mem[3029] = 4'b0110;
	mem[3030] = 4'b0110;
	mem[3031] = 4'b0110;
	mem[3032] = 4'b0110;
	mem[3033] = 4'b0110;
	mem[3034] = 4'b0110;
	mem[3035] = 4'b0110;
	mem[3036] = 4'b0110;
	mem[3037] = 4'b0110;
	mem[3038] = 4'b0110;
	mem[3039] = 4'b0110;
	mem[3040] = 4'b0110;
	mem[3041] = 4'b0110;
	mem[3042] = 4'b0110;
	mem[3043] = 4'b0110;
	mem[3044] = 4'b0110;
	mem[3045] = 4'b0110;
	mem[3046] = 4'b0110;
	mem[3047] = 4'b0110;
	mem[3048] = 4'b0111;
	mem[3049] = 4'b0111;
	mem[3050] = 4'b0111;
	mem[3051] = 4'b0111;
	mem[3052] = 4'b0111;
	mem[3053] = 4'b0110;
	mem[3054] = 4'b0110;
	mem[3055] = 4'b0110;
	mem[3056] = 4'b0110;
	mem[3057] = 4'b0110;
	mem[3058] = 4'b0110;
	mem[3059] = 4'b0110;
	mem[3060] = 4'b0110;
	mem[3061] = 4'b0111;
	mem[3062] = 4'b1000;
	mem[3063] = 4'b0111;
	mem[3064] = 4'b0000;
	mem[3065] = 4'b0000;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b0111;
	mem[3076] = 4'b1100;
	mem[3077] = 4'b1101;
	mem[3078] = 4'b1101;
	mem[3079] = 4'b1101;
	mem[3080] = 4'b1101;
	mem[3081] = 4'b1101;
	mem[3082] = 4'b1101;
	mem[3083] = 4'b1101;
	mem[3084] = 4'b1101;
	mem[3085] = 4'b1101;
	mem[3086] = 4'b1101;
	mem[3087] = 4'b1101;
	mem[3088] = 4'b1101;
	mem[3089] = 4'b1101;
	mem[3090] = 4'b1101;
	mem[3091] = 4'b1101;
	mem[3092] = 4'b1111;
	mem[3093] = 4'b1111;
	mem[3094] = 4'b1111;
	mem[3095] = 4'b1111;
	mem[3096] = 4'b1111;
	mem[3097] = 4'b1111;
	mem[3098] = 4'b1111;
	mem[3099] = 4'b1111;
	mem[3100] = 4'b1111;
	mem[3101] = 4'b1111;
	mem[3102] = 4'b1111;
	mem[3103] = 4'b1111;
	mem[3104] = 4'b1111;
	mem[3105] = 4'b1111;
	mem[3106] = 4'b1111;
	mem[3107] = 4'b1111;
	mem[3108] = 4'b1111;
	mem[3109] = 4'b1111;
	mem[3110] = 4'b1111;
	mem[3111] = 4'b1111;
	mem[3112] = 4'b1111;
	mem[3113] = 4'b1111;
	mem[3114] = 4'b1111;
	mem[3115] = 4'b1111;
	mem[3116] = 4'b1111;
	mem[3117] = 4'b1111;
	mem[3118] = 4'b1111;
	mem[3119] = 4'b1111;
	mem[3120] = 4'b1110;
	mem[3121] = 4'b1101;
	mem[3122] = 4'b1111;
	mem[3123] = 4'b1111;
	mem[3124] = 4'b1110;
	mem[3125] = 4'b1110;
	mem[3126] = 4'b1110;
	mem[3127] = 4'b1101;
	mem[3128] = 4'b1101;
	mem[3129] = 4'b1111;
	mem[3130] = 4'b1111;
	mem[3131] = 4'b1111;
	mem[3132] = 4'b1111;
	mem[3133] = 4'b1111;
	mem[3134] = 4'b1111;
	mem[3135] = 4'b1111;
	mem[3136] = 4'b1111;
	mem[3137] = 4'b1111;
	mem[3138] = 4'b1111;
	mem[3139] = 4'b1111;
	mem[3140] = 4'b1111;
	mem[3141] = 4'b1111;
	mem[3142] = 4'b1111;
	mem[3143] = 4'b1000;
	mem[3144] = 4'b0110;
	mem[3145] = 4'b0110;
	mem[3146] = 4'b0110;
	mem[3147] = 4'b0110;
	mem[3148] = 4'b0110;
	mem[3149] = 4'b0110;
	mem[3150] = 4'b0110;
	mem[3151] = 4'b0110;
	mem[3152] = 4'b0110;
	mem[3153] = 4'b0110;
	mem[3154] = 4'b0110;
	mem[3155] = 4'b0110;
	mem[3156] = 4'b0110;
	mem[3157] = 4'b0110;
	mem[3158] = 4'b0110;
	mem[3159] = 4'b0110;
	mem[3160] = 4'b0110;
	mem[3161] = 4'b0110;
	mem[3162] = 4'b0110;
	mem[3163] = 4'b0110;
	mem[3164] = 4'b0110;
	mem[3165] = 4'b0110;
	mem[3166] = 4'b0110;
	mem[3167] = 4'b0110;
	mem[3168] = 4'b0110;
	mem[3169] = 4'b0110;
	mem[3170] = 4'b0110;
	mem[3171] = 4'b0110;
	mem[3172] = 4'b0110;
	mem[3173] = 4'b0110;
	mem[3174] = 4'b0110;
	mem[3175] = 4'b0110;
	mem[3176] = 4'b0110;
	mem[3177] = 4'b0111;
	mem[3178] = 4'b0111;
	mem[3179] = 4'b0111;
	mem[3180] = 4'b0111;
	mem[3181] = 4'b0111;
	mem[3182] = 4'b0111;
	mem[3183] = 4'b0110;
	mem[3184] = 4'b0110;
	mem[3185] = 4'b0110;
	mem[3186] = 4'b0110;
	mem[3187] = 4'b0111;
	mem[3188] = 4'b1000;
	mem[3189] = 4'b1000;
	mem[3190] = 4'b0111;
	mem[3191] = 4'b0111;
	mem[3192] = 4'b0000;
	mem[3193] = 4'b0000;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b0111;
	mem[3204] = 4'b1100;
	mem[3205] = 4'b1101;
	mem[3206] = 4'b1101;
	mem[3207] = 4'b1101;
	mem[3208] = 4'b1101;
	mem[3209] = 4'b1101;
	mem[3210] = 4'b1101;
	mem[3211] = 4'b1101;
	mem[3212] = 4'b1101;
	mem[3213] = 4'b1101;
	mem[3214] = 4'b1101;
	mem[3215] = 4'b1101;
	mem[3216] = 4'b1101;
	mem[3217] = 4'b1101;
	mem[3218] = 4'b1101;
	mem[3219] = 4'b1101;
	mem[3220] = 4'b1111;
	mem[3221] = 4'b1111;
	mem[3222] = 4'b1111;
	mem[3223] = 4'b1111;
	mem[3224] = 4'b1111;
	mem[3225] = 4'b1111;
	mem[3226] = 4'b1111;
	mem[3227] = 4'b1111;
	mem[3228] = 4'b1111;
	mem[3229] = 4'b1111;
	mem[3230] = 4'b1111;
	mem[3231] = 4'b1111;
	mem[3232] = 4'b1111;
	mem[3233] = 4'b1111;
	mem[3234] = 4'b1111;
	mem[3235] = 4'b1111;
	mem[3236] = 4'b1111;
	mem[3237] = 4'b1111;
	mem[3238] = 4'b1111;
	mem[3239] = 4'b1111;
	mem[3240] = 4'b1111;
	mem[3241] = 4'b1111;
	mem[3242] = 4'b1111;
	mem[3243] = 4'b1111;
	mem[3244] = 4'b1111;
	mem[3245] = 4'b1111;
	mem[3246] = 4'b1111;
	mem[3247] = 4'b1111;
	mem[3248] = 4'b1111;
	mem[3249] = 4'b1110;
	mem[3250] = 4'b1111;
	mem[3251] = 4'b1111;
	mem[3252] = 4'b1101;
	mem[3253] = 4'b1111;
	mem[3254] = 4'b1111;
	mem[3255] = 4'b1110;
	mem[3256] = 4'b1101;
	mem[3257] = 4'b1101;
	mem[3258] = 4'b1110;
	mem[3259] = 4'b1111;
	mem[3260] = 4'b1111;
	mem[3261] = 4'b1111;
	mem[3262] = 4'b1111;
	mem[3263] = 4'b1111;
	mem[3264] = 4'b1111;
	mem[3265] = 4'b1111;
	mem[3266] = 4'b1111;
	mem[3267] = 4'b1111;
	mem[3268] = 4'b1111;
	mem[3269] = 4'b1111;
	mem[3270] = 4'b1111;
	mem[3271] = 4'b1000;
	mem[3272] = 4'b0110;
	mem[3273] = 4'b0110;
	mem[3274] = 4'b0110;
	mem[3275] = 4'b0110;
	mem[3276] = 4'b0110;
	mem[3277] = 4'b0110;
	mem[3278] = 4'b0110;
	mem[3279] = 4'b0110;
	mem[3280] = 4'b0110;
	mem[3281] = 4'b0110;
	mem[3282] = 4'b0110;
	mem[3283] = 4'b0110;
	mem[3284] = 4'b0110;
	mem[3285] = 4'b0110;
	mem[3286] = 4'b0110;
	mem[3287] = 4'b0110;
	mem[3288] = 4'b0110;
	mem[3289] = 4'b0110;
	mem[3290] = 4'b0110;
	mem[3291] = 4'b0110;
	mem[3292] = 4'b0110;
	mem[3293] = 4'b0110;
	mem[3294] = 4'b0110;
	mem[3295] = 4'b0110;
	mem[3296] = 4'b0110;
	mem[3297] = 4'b0110;
	mem[3298] = 4'b0111;
	mem[3299] = 4'b0111;
	mem[3300] = 4'b0110;
	mem[3301] = 4'b0110;
	mem[3302] = 4'b0110;
	mem[3303] = 4'b0110;
	mem[3304] = 4'b0110;
	mem[3305] = 4'b0110;
	mem[3306] = 4'b0111;
	mem[3307] = 4'b0111;
	mem[3308] = 4'b0111;
	mem[3309] = 4'b0111;
	mem[3310] = 4'b0111;
	mem[3311] = 4'b0111;
	mem[3312] = 4'b0111;
	mem[3313] = 4'b1000;
	mem[3314] = 4'b1000;
	mem[3315] = 4'b1000;
	mem[3316] = 4'b0111;
	mem[3317] = 4'b0111;
	mem[3318] = 4'b0111;
	mem[3319] = 4'b0111;
	mem[3320] = 4'b0000;
	mem[3321] = 4'b0000;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b0111;
	mem[3332] = 4'b1100;
	mem[3333] = 4'b1101;
	mem[3334] = 4'b1101;
	mem[3335] = 4'b1101;
	mem[3336] = 4'b1101;
	mem[3337] = 4'b1101;
	mem[3338] = 4'b1101;
	mem[3339] = 4'b1101;
	mem[3340] = 4'b1101;
	mem[3341] = 4'b1101;
	mem[3342] = 4'b1101;
	mem[3343] = 4'b1101;
	mem[3344] = 4'b1101;
	mem[3345] = 4'b1101;
	mem[3346] = 4'b1101;
	mem[3347] = 4'b1101;
	mem[3348] = 4'b1111;
	mem[3349] = 4'b1111;
	mem[3350] = 4'b1111;
	mem[3351] = 4'b1111;
	mem[3352] = 4'b1111;
	mem[3353] = 4'b1111;
	mem[3354] = 4'b1111;
	mem[3355] = 4'b1111;
	mem[3356] = 4'b1111;
	mem[3357] = 4'b1111;
	mem[3358] = 4'b1111;
	mem[3359] = 4'b1111;
	mem[3360] = 4'b1111;
	mem[3361] = 4'b1111;
	mem[3362] = 4'b1111;
	mem[3363] = 4'b1111;
	mem[3364] = 4'b1111;
	mem[3365] = 4'b1111;
	mem[3366] = 4'b1111;
	mem[3367] = 4'b1111;
	mem[3368] = 4'b1111;
	mem[3369] = 4'b1111;
	mem[3370] = 4'b1111;
	mem[3371] = 4'b1111;
	mem[3372] = 4'b1111;
	mem[3373] = 4'b1111;
	mem[3374] = 4'b1111;
	mem[3375] = 4'b1111;
	mem[3376] = 4'b1111;
	mem[3377] = 4'b1111;
	mem[3378] = 4'b1111;
	mem[3379] = 4'b1110;
	mem[3380] = 4'b1110;
	mem[3381] = 4'b1111;
	mem[3382] = 4'b1111;
	mem[3383] = 4'b1110;
	mem[3384] = 4'b1110;
	mem[3385] = 4'b1110;
	mem[3386] = 4'b1111;
	mem[3387] = 4'b1111;
	mem[3388] = 4'b1111;
	mem[3389] = 4'b1111;
	mem[3390] = 4'b1111;
	mem[3391] = 4'b1111;
	mem[3392] = 4'b1111;
	mem[3393] = 4'b1111;
	mem[3394] = 4'b1111;
	mem[3395] = 4'b1111;
	mem[3396] = 4'b1111;
	mem[3397] = 4'b1111;
	mem[3398] = 4'b1111;
	mem[3399] = 4'b1000;
	mem[3400] = 4'b0110;
	mem[3401] = 4'b0110;
	mem[3402] = 4'b0110;
	mem[3403] = 4'b0110;
	mem[3404] = 4'b0110;
	mem[3405] = 4'b0110;
	mem[3406] = 4'b0110;
	mem[3407] = 4'b0110;
	mem[3408] = 4'b0110;
	mem[3409] = 4'b0110;
	mem[3410] = 4'b0110;
	mem[3411] = 4'b0110;
	mem[3412] = 4'b0110;
	mem[3413] = 4'b0110;
	mem[3414] = 4'b0110;
	mem[3415] = 4'b0110;
	mem[3416] = 4'b0110;
	mem[3417] = 4'b0110;
	mem[3418] = 4'b0110;
	mem[3419] = 4'b0110;
	mem[3420] = 4'b0110;
	mem[3421] = 4'b0110;
	mem[3422] = 4'b0110;
	mem[3423] = 4'b0110;
	mem[3424] = 4'b0110;
	mem[3425] = 4'b0111;
	mem[3426] = 4'b0111;
	mem[3427] = 4'b0111;
	mem[3428] = 4'b0111;
	mem[3429] = 4'b0110;
	mem[3430] = 4'b0110;
	mem[3431] = 4'b0110;
	mem[3432] = 4'b0110;
	mem[3433] = 4'b0110;
	mem[3434] = 4'b0111;
	mem[3435] = 4'b0111;
	mem[3436] = 4'b0111;
	mem[3437] = 4'b0111;
	mem[3438] = 4'b0111;
	mem[3439] = 4'b0111;
	mem[3440] = 4'b0111;
	mem[3441] = 4'b0111;
	mem[3442] = 4'b0111;
	mem[3443] = 4'b0111;
	mem[3444] = 4'b0111;
	mem[3445] = 4'b0111;
	mem[3446] = 4'b0111;
	mem[3447] = 4'b0111;
	mem[3448] = 4'b0000;
	mem[3449] = 4'b0000;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b0111;
	mem[3460] = 4'b1100;
	mem[3461] = 4'b1101;
	mem[3462] = 4'b1101;
	mem[3463] = 4'b1101;
	mem[3464] = 4'b1101;
	mem[3465] = 4'b1101;
	mem[3466] = 4'b1101;
	mem[3467] = 4'b1101;
	mem[3468] = 4'b1101;
	mem[3469] = 4'b1101;
	mem[3470] = 4'b1101;
	mem[3471] = 4'b1101;
	mem[3472] = 4'b1101;
	mem[3473] = 4'b1101;
	mem[3474] = 4'b1101;
	mem[3475] = 4'b1101;
	mem[3476] = 4'b1111;
	mem[3477] = 4'b1111;
	mem[3478] = 4'b1111;
	mem[3479] = 4'b1111;
	mem[3480] = 4'b1111;
	mem[3481] = 4'b1111;
	mem[3482] = 4'b1111;
	mem[3483] = 4'b1111;
	mem[3484] = 4'b1111;
	mem[3485] = 4'b1111;
	mem[3486] = 4'b1111;
	mem[3487] = 4'b1111;
	mem[3488] = 4'b1111;
	mem[3489] = 4'b1111;
	mem[3490] = 4'b1111;
	mem[3491] = 4'b1111;
	mem[3492] = 4'b1111;
	mem[3493] = 4'b1111;
	mem[3494] = 4'b1111;
	mem[3495] = 4'b1111;
	mem[3496] = 4'b1111;
	mem[3497] = 4'b1111;
	mem[3498] = 4'b1111;
	mem[3499] = 4'b1111;
	mem[3500] = 4'b1111;
	mem[3501] = 4'b1111;
	mem[3502] = 4'b1111;
	mem[3503] = 4'b1111;
	mem[3504] = 4'b1111;
	mem[3505] = 4'b1111;
	mem[3506] = 4'b1111;
	mem[3507] = 4'b1101;
	mem[3508] = 4'b1110;
	mem[3509] = 4'b1111;
	mem[3510] = 4'b1111;
	mem[3511] = 4'b1101;
	mem[3512] = 4'b1111;
	mem[3513] = 4'b1111;
	mem[3514] = 4'b1111;
	mem[3515] = 4'b1111;
	mem[3516] = 4'b1111;
	mem[3517] = 4'b1111;
	mem[3518] = 4'b1111;
	mem[3519] = 4'b1111;
	mem[3520] = 4'b1111;
	mem[3521] = 4'b1111;
	mem[3522] = 4'b1111;
	mem[3523] = 4'b1111;
	mem[3524] = 4'b1111;
	mem[3525] = 4'b1111;
	mem[3526] = 4'b1111;
	mem[3527] = 4'b1000;
	mem[3528] = 4'b0110;
	mem[3529] = 4'b0110;
	mem[3530] = 4'b0110;
	mem[3531] = 4'b0110;
	mem[3532] = 4'b0110;
	mem[3533] = 4'b0110;
	mem[3534] = 4'b0110;
	mem[3535] = 4'b0110;
	mem[3536] = 4'b0110;
	mem[3537] = 4'b0110;
	mem[3538] = 4'b0110;
	mem[3539] = 4'b0110;
	mem[3540] = 4'b0110;
	mem[3541] = 4'b0110;
	mem[3542] = 4'b0110;
	mem[3543] = 4'b0110;
	mem[3544] = 4'b0110;
	mem[3545] = 4'b0110;
	mem[3546] = 4'b0110;
	mem[3547] = 4'b0110;
	mem[3548] = 4'b0110;
	mem[3549] = 4'b0110;
	mem[3550] = 4'b0111;
	mem[3551] = 4'b0110;
	mem[3552] = 4'b0111;
	mem[3553] = 4'b0111;
	mem[3554] = 4'b0111;
	mem[3555] = 4'b0111;
	mem[3556] = 4'b0111;
	mem[3557] = 4'b0111;
	mem[3558] = 4'b0110;
	mem[3559] = 4'b0110;
	mem[3560] = 4'b0110;
	mem[3561] = 4'b0110;
	mem[3562] = 4'b0110;
	mem[3563] = 4'b0111;
	mem[3564] = 4'b0111;
	mem[3565] = 4'b0111;
	mem[3566] = 4'b0111;
	mem[3567] = 4'b0111;
	mem[3568] = 4'b0111;
	mem[3569] = 4'b0111;
	mem[3570] = 4'b0111;
	mem[3571] = 4'b0111;
	mem[3572] = 4'b0111;
	mem[3573] = 4'b0111;
	mem[3574] = 4'b0111;
	mem[3575] = 4'b0111;
	mem[3576] = 4'b0000;
	mem[3577] = 4'b0000;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b0111;
	mem[3588] = 4'b1100;
	mem[3589] = 4'b1101;
	mem[3590] = 4'b1101;
	mem[3591] = 4'b1101;
	mem[3592] = 4'b1101;
	mem[3593] = 4'b1101;
	mem[3594] = 4'b1101;
	mem[3595] = 4'b1101;
	mem[3596] = 4'b1101;
	mem[3597] = 4'b1101;
	mem[3598] = 4'b1101;
	mem[3599] = 4'b1101;
	mem[3600] = 4'b1101;
	mem[3601] = 4'b1101;
	mem[3602] = 4'b1101;
	mem[3603] = 4'b1101;
	mem[3604] = 4'b1111;
	mem[3605] = 4'b1111;
	mem[3606] = 4'b1111;
	mem[3607] = 4'b1111;
	mem[3608] = 4'b1111;
	mem[3609] = 4'b1111;
	mem[3610] = 4'b1111;
	mem[3611] = 4'b1111;
	mem[3612] = 4'b1111;
	mem[3613] = 4'b1111;
	mem[3614] = 4'b1111;
	mem[3615] = 4'b1111;
	mem[3616] = 4'b1111;
	mem[3617] = 4'b1111;
	mem[3618] = 4'b1111;
	mem[3619] = 4'b1111;
	mem[3620] = 4'b1111;
	mem[3621] = 4'b1111;
	mem[3622] = 4'b1111;
	mem[3623] = 4'b1101;
	mem[3624] = 4'b1110;
	mem[3625] = 4'b1111;
	mem[3626] = 4'b1111;
	mem[3627] = 4'b1111;
	mem[3628] = 4'b1111;
	mem[3629] = 4'b1111;
	mem[3630] = 4'b1111;
	mem[3631] = 4'b1111;
	mem[3632] = 4'b1111;
	mem[3633] = 4'b1111;
	mem[3634] = 4'b1111;
	mem[3635] = 4'b1101;
	mem[3636] = 4'b1101;
	mem[3637] = 4'b1101;
	mem[3638] = 4'b1101;
	mem[3639] = 4'b1110;
	mem[3640] = 4'b1111;
	mem[3641] = 4'b1111;
	mem[3642] = 4'b1111;
	mem[3643] = 4'b1111;
	mem[3644] = 4'b1111;
	mem[3645] = 4'b1111;
	mem[3646] = 4'b1111;
	mem[3647] = 4'b1111;
	mem[3648] = 4'b1111;
	mem[3649] = 4'b1111;
	mem[3650] = 4'b1111;
	mem[3651] = 4'b1111;
	mem[3652] = 4'b1111;
	mem[3653] = 4'b1111;
	mem[3654] = 4'b1111;
	mem[3655] = 4'b1000;
	mem[3656] = 4'b0110;
	mem[3657] = 4'b0110;
	mem[3658] = 4'b0110;
	mem[3659] = 4'b0110;
	mem[3660] = 4'b0110;
	mem[3661] = 4'b0110;
	mem[3662] = 4'b0110;
	mem[3663] = 4'b0110;
	mem[3664] = 4'b0110;
	mem[3665] = 4'b0110;
	mem[3666] = 4'b0110;
	mem[3667] = 4'b0110;
	mem[3668] = 4'b0110;
	mem[3669] = 4'b0110;
	mem[3670] = 4'b0110;
	mem[3671] = 4'b0110;
	mem[3672] = 4'b0110;
	mem[3673] = 4'b0110;
	mem[3674] = 4'b0110;
	mem[3675] = 4'b0110;
	mem[3676] = 4'b0110;
	mem[3677] = 4'b0110;
	mem[3678] = 4'b0110;
	mem[3679] = 4'b0110;
	mem[3680] = 4'b0111;
	mem[3681] = 4'b0111;
	mem[3682] = 4'b0111;
	mem[3683] = 4'b0111;
	mem[3684] = 4'b0111;
	mem[3685] = 4'b0111;
	mem[3686] = 4'b0111;
	mem[3687] = 4'b0111;
	mem[3688] = 4'b0110;
	mem[3689] = 4'b0110;
	mem[3690] = 4'b0110;
	mem[3691] = 4'b0110;
	mem[3692] = 4'b0111;
	mem[3693] = 4'b0111;
	mem[3694] = 4'b0111;
	mem[3695] = 4'b0111;
	mem[3696] = 4'b0111;
	mem[3697] = 4'b0111;
	mem[3698] = 4'b0111;
	mem[3699] = 4'b0111;
	mem[3700] = 4'b0111;
	mem[3701] = 4'b0111;
	mem[3702] = 4'b0111;
	mem[3703] = 4'b0111;
	mem[3704] = 4'b0000;
	mem[3705] = 4'b0000;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b0111;
	mem[3716] = 4'b1100;
	mem[3717] = 4'b1101;
	mem[3718] = 4'b1101;
	mem[3719] = 4'b1101;
	mem[3720] = 4'b1101;
	mem[3721] = 4'b1101;
	mem[3722] = 4'b1101;
	mem[3723] = 4'b1101;
	mem[3724] = 4'b1101;
	mem[3725] = 4'b1101;
	mem[3726] = 4'b1101;
	mem[3727] = 4'b1101;
	mem[3728] = 4'b1101;
	mem[3729] = 4'b1101;
	mem[3730] = 4'b1101;
	mem[3731] = 4'b1101;
	mem[3732] = 4'b1111;
	mem[3733] = 4'b1111;
	mem[3734] = 4'b1111;
	mem[3735] = 4'b1111;
	mem[3736] = 4'b1111;
	mem[3737] = 4'b1111;
	mem[3738] = 4'b1111;
	mem[3739] = 4'b1111;
	mem[3740] = 4'b1111;
	mem[3741] = 4'b1111;
	mem[3742] = 4'b1111;
	mem[3743] = 4'b1111;
	mem[3744] = 4'b1111;
	mem[3745] = 4'b1111;
	mem[3746] = 4'b1111;
	mem[3747] = 4'b1111;
	mem[3748] = 4'b1111;
	mem[3749] = 4'b1111;
	mem[3750] = 4'b1110;
	mem[3751] = 4'b1101;
	mem[3752] = 4'b1101;
	mem[3753] = 4'b1110;
	mem[3754] = 4'b1111;
	mem[3755] = 4'b1111;
	mem[3756] = 4'b1111;
	mem[3757] = 4'b1111;
	mem[3758] = 4'b1111;
	mem[3759] = 4'b1111;
	mem[3760] = 4'b1111;
	mem[3761] = 4'b1111;
	mem[3762] = 4'b1111;
	mem[3763] = 4'b1111;
	mem[3764] = 4'b1110;
	mem[3765] = 4'b1101;
	mem[3766] = 4'b1110;
	mem[3767] = 4'b1111;
	mem[3768] = 4'b1111;
	mem[3769] = 4'b1111;
	mem[3770] = 4'b1111;
	mem[3771] = 4'b1111;
	mem[3772] = 4'b1111;
	mem[3773] = 4'b1111;
	mem[3774] = 4'b1111;
	mem[3775] = 4'b1111;
	mem[3776] = 4'b1111;
	mem[3777] = 4'b1111;
	mem[3778] = 4'b1111;
	mem[3779] = 4'b1111;
	mem[3780] = 4'b1111;
	mem[3781] = 4'b1111;
	mem[3782] = 4'b1111;
	mem[3783] = 4'b1000;
	mem[3784] = 4'b0110;
	mem[3785] = 4'b0110;
	mem[3786] = 4'b0110;
	mem[3787] = 4'b0110;
	mem[3788] = 4'b0110;
	mem[3789] = 4'b0110;
	mem[3790] = 4'b0110;
	mem[3791] = 4'b0110;
	mem[3792] = 4'b0110;
	mem[3793] = 4'b0110;
	mem[3794] = 4'b0110;
	mem[3795] = 4'b0110;
	mem[3796] = 4'b0110;
	mem[3797] = 4'b0110;
	mem[3798] = 4'b0110;
	mem[3799] = 4'b0110;
	mem[3800] = 4'b0110;
	mem[3801] = 4'b0111;
	mem[3802] = 4'b0111;
	mem[3803] = 4'b0110;
	mem[3804] = 4'b0110;
	mem[3805] = 4'b0110;
	mem[3806] = 4'b0110;
	mem[3807] = 4'b0110;
	mem[3808] = 4'b0111;
	mem[3809] = 4'b0111;
	mem[3810] = 4'b0111;
	mem[3811] = 4'b0111;
	mem[3812] = 4'b0111;
	mem[3813] = 4'b0111;
	mem[3814] = 4'b0111;
	mem[3815] = 4'b0111;
	mem[3816] = 4'b0111;
	mem[3817] = 4'b0110;
	mem[3818] = 4'b0110;
	mem[3819] = 4'b0110;
	mem[3820] = 4'b0110;
	mem[3821] = 4'b0111;
	mem[3822] = 4'b0111;
	mem[3823] = 4'b0111;
	mem[3824] = 4'b0111;
	mem[3825] = 4'b0111;
	mem[3826] = 4'b0111;
	mem[3827] = 4'b0111;
	mem[3828] = 4'b0111;
	mem[3829] = 4'b0111;
	mem[3830] = 4'b0111;
	mem[3831] = 4'b0111;
	mem[3832] = 4'b0000;
	mem[3833] = 4'b0000;
	mem[3834] = 4'b0000;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b0111;
	mem[3844] = 4'b1100;
	mem[3845] = 4'b1101;
	mem[3846] = 4'b1101;
	mem[3847] = 4'b1101;
	mem[3848] = 4'b1101;
	mem[3849] = 4'b1101;
	mem[3850] = 4'b1101;
	mem[3851] = 4'b1101;
	mem[3852] = 4'b1101;
	mem[3853] = 4'b1101;
	mem[3854] = 4'b1101;
	mem[3855] = 4'b1101;
	mem[3856] = 4'b1101;
	mem[3857] = 4'b1101;
	mem[3858] = 4'b1101;
	mem[3859] = 4'b1101;
	mem[3860] = 4'b1111;
	mem[3861] = 4'b1111;
	mem[3862] = 4'b1111;
	mem[3863] = 4'b1111;
	mem[3864] = 4'b1111;
	mem[3865] = 4'b1111;
	mem[3866] = 4'b1111;
	mem[3867] = 4'b1111;
	mem[3868] = 4'b1111;
	mem[3869] = 4'b1111;
	mem[3870] = 4'b1111;
	mem[3871] = 4'b1111;
	mem[3872] = 4'b1111;
	mem[3873] = 4'b1111;
	mem[3874] = 4'b1111;
	mem[3875] = 4'b1111;
	mem[3876] = 4'b1111;
	mem[3877] = 4'b1111;
	mem[3878] = 4'b1111;
	mem[3879] = 4'b1110;
	mem[3880] = 4'b1101;
	mem[3881] = 4'b1101;
	mem[3882] = 4'b1110;
	mem[3883] = 4'b1111;
	mem[3884] = 4'b1111;
	mem[3885] = 4'b1111;
	mem[3886] = 4'b1111;
	mem[3887] = 4'b1111;
	mem[3888] = 4'b1111;
	mem[3889] = 4'b1111;
	mem[3890] = 4'b1111;
	mem[3891] = 4'b1111;
	mem[3892] = 4'b1111;
	mem[3893] = 4'b1111;
	mem[3894] = 4'b1111;
	mem[3895] = 4'b1111;
	mem[3896] = 4'b1111;
	mem[3897] = 4'b1111;
	mem[3898] = 4'b1111;
	mem[3899] = 4'b1111;
	mem[3900] = 4'b1111;
	mem[3901] = 4'b1111;
	mem[3902] = 4'b1111;
	mem[3903] = 4'b1111;
	mem[3904] = 4'b1111;
	mem[3905] = 4'b1111;
	mem[3906] = 4'b1111;
	mem[3907] = 4'b1111;
	mem[3908] = 4'b1111;
	mem[3909] = 4'b1111;
	mem[3910] = 4'b1111;
	mem[3911] = 4'b1001;
	mem[3912] = 4'b0110;
	mem[3913] = 4'b0110;
	mem[3914] = 4'b0110;
	mem[3915] = 4'b0110;
	mem[3916] = 4'b0110;
	mem[3917] = 4'b0110;
	mem[3918] = 4'b0110;
	mem[3919] = 4'b0110;
	mem[3920] = 4'b0110;
	mem[3921] = 4'b0110;
	mem[3922] = 4'b0110;
	mem[3923] = 4'b0110;
	mem[3924] = 4'b0110;
	mem[3925] = 4'b0110;
	mem[3926] = 4'b0110;
	mem[3927] = 4'b0111;
	mem[3928] = 4'b0111;
	mem[3929] = 4'b0111;
	mem[3930] = 4'b0111;
	mem[3931] = 4'b0111;
	mem[3932] = 4'b0110;
	mem[3933] = 4'b0110;
	mem[3934] = 4'b0110;
	mem[3935] = 4'b0110;
	mem[3936] = 4'b0110;
	mem[3937] = 4'b0111;
	mem[3938] = 4'b0111;
	mem[3939] = 4'b0111;
	mem[3940] = 4'b0111;
	mem[3941] = 4'b0111;
	mem[3942] = 4'b0111;
	mem[3943] = 4'b0111;
	mem[3944] = 4'b0111;
	mem[3945] = 4'b0111;
	mem[3946] = 4'b0110;
	mem[3947] = 4'b0110;
	mem[3948] = 4'b0110;
	mem[3949] = 4'b0110;
	mem[3950] = 4'b0111;
	mem[3951] = 4'b0111;
	mem[3952] = 4'b0111;
	mem[3953] = 4'b0111;
	mem[3954] = 4'b0111;
	mem[3955] = 4'b0111;
	mem[3956] = 4'b0111;
	mem[3957] = 4'b0111;
	mem[3958] = 4'b0111;
	mem[3959] = 4'b0111;
	mem[3960] = 4'b0000;
	mem[3961] = 4'b0000;
	mem[3962] = 4'b0000;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b0111;
	mem[3972] = 4'b1100;
	mem[3973] = 4'b1101;
	mem[3974] = 4'b1101;
	mem[3975] = 4'b1101;
	mem[3976] = 4'b1101;
	mem[3977] = 4'b1101;
	mem[3978] = 4'b1101;
	mem[3979] = 4'b1101;
	mem[3980] = 4'b1101;
	mem[3981] = 4'b1101;
	mem[3982] = 4'b1101;
	mem[3983] = 4'b1101;
	mem[3984] = 4'b1101;
	mem[3985] = 4'b1101;
	mem[3986] = 4'b1101;
	mem[3987] = 4'b1101;
	mem[3988] = 4'b1111;
	mem[3989] = 4'b1111;
	mem[3990] = 4'b1111;
	mem[3991] = 4'b1111;
	mem[3992] = 4'b1111;
	mem[3993] = 4'b1111;
	mem[3994] = 4'b1111;
	mem[3995] = 4'b1111;
	mem[3996] = 4'b1111;
	mem[3997] = 4'b1111;
	mem[3998] = 4'b1111;
	mem[3999] = 4'b1111;
	mem[4000] = 4'b1111;
	mem[4001] = 4'b1111;
	mem[4002] = 4'b1111;
	mem[4003] = 4'b1111;
	mem[4004] = 4'b1111;
	mem[4005] = 4'b1111;
	mem[4006] = 4'b1111;
	mem[4007] = 4'b1111;
	mem[4008] = 4'b1110;
	mem[4009] = 4'b1101;
	mem[4010] = 4'b1101;
	mem[4011] = 4'b1110;
	mem[4012] = 4'b1111;
	mem[4013] = 4'b1111;
	mem[4014] = 4'b1111;
	mem[4015] = 4'b1111;
	mem[4016] = 4'b1111;
	mem[4017] = 4'b1111;
	mem[4018] = 4'b1101;
	mem[4019] = 4'b1101;
	mem[4020] = 4'b1111;
	mem[4021] = 4'b1111;
	mem[4022] = 4'b1111;
	mem[4023] = 4'b1111;
	mem[4024] = 4'b1111;
	mem[4025] = 4'b1111;
	mem[4026] = 4'b1111;
	mem[4027] = 4'b1111;
	mem[4028] = 4'b1111;
	mem[4029] = 4'b1111;
	mem[4030] = 4'b1111;
	mem[4031] = 4'b1111;
	mem[4032] = 4'b1111;
	mem[4033] = 4'b1111;
	mem[4034] = 4'b1111;
	mem[4035] = 4'b1111;
	mem[4036] = 4'b1111;
	mem[4037] = 4'b1111;
	mem[4038] = 4'b1111;
	mem[4039] = 4'b1001;
	mem[4040] = 4'b0110;
	mem[4041] = 4'b0110;
	mem[4042] = 4'b0110;
	mem[4043] = 4'b0110;
	mem[4044] = 4'b0110;
	mem[4045] = 4'b0110;
	mem[4046] = 4'b0110;
	mem[4047] = 4'b0110;
	mem[4048] = 4'b0110;
	mem[4049] = 4'b0110;
	mem[4050] = 4'b0110;
	mem[4051] = 4'b0110;
	mem[4052] = 4'b0110;
	mem[4053] = 4'b0111;
	mem[4054] = 4'b0111;
	mem[4055] = 4'b0111;
	mem[4056] = 4'b0111;
	mem[4057] = 4'b0111;
	mem[4058] = 4'b0111;
	mem[4059] = 4'b0111;
	mem[4060] = 4'b0111;
	mem[4061] = 4'b0110;
	mem[4062] = 4'b0110;
	mem[4063] = 4'b0110;
	mem[4064] = 4'b0110;
	mem[4065] = 4'b0110;
	mem[4066] = 4'b0111;
	mem[4067] = 4'b0111;
	mem[4068] = 4'b0111;
	mem[4069] = 4'b0111;
	mem[4070] = 4'b0111;
	mem[4071] = 4'b0111;
	mem[4072] = 4'b0111;
	mem[4073] = 4'b0111;
	mem[4074] = 4'b0111;
	mem[4075] = 4'b0110;
	mem[4076] = 4'b0110;
	mem[4077] = 4'b0111;
	mem[4078] = 4'b1000;
	mem[4079] = 4'b0111;
	mem[4080] = 4'b0111;
	mem[4081] = 4'b0111;
	mem[4082] = 4'b0111;
	mem[4083] = 4'b0111;
	mem[4084] = 4'b0111;
	mem[4085] = 4'b0111;
	mem[4086] = 4'b0111;
	mem[4087] = 4'b0111;
	mem[4088] = 4'b0000;
	mem[4089] = 4'b0000;
	mem[4090] = 4'b0000;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_1g (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0111;
	mem[4] = 4'b1100;
	mem[5] = 4'b1101;
	mem[6] = 4'b1101;
	mem[7] = 4'b1101;
	mem[8] = 4'b1101;
	mem[9] = 4'b1101;
	mem[10] = 4'b1101;
	mem[11] = 4'b1101;
	mem[12] = 4'b1101;
	mem[13] = 4'b1101;
	mem[14] = 4'b1101;
	mem[15] = 4'b1101;
	mem[16] = 4'b1101;
	mem[17] = 4'b1101;
	mem[18] = 4'b1101;
	mem[19] = 4'b1101;
	mem[20] = 4'b1111;
	mem[21] = 4'b1111;
	mem[22] = 4'b1111;
	mem[23] = 4'b1111;
	mem[24] = 4'b1111;
	mem[25] = 4'b1111;
	mem[26] = 4'b1111;
	mem[27] = 4'b1111;
	mem[28] = 4'b1111;
	mem[29] = 4'b1111;
	mem[30] = 4'b1111;
	mem[31] = 4'b1111;
	mem[32] = 4'b1111;
	mem[33] = 4'b1111;
	mem[34] = 4'b1111;
	mem[35] = 4'b1111;
	mem[36] = 4'b1111;
	mem[37] = 4'b1111;
	mem[38] = 4'b1111;
	mem[39] = 4'b1111;
	mem[40] = 4'b1111;
	mem[41] = 4'b1110;
	mem[42] = 4'b1101;
	mem[43] = 4'b1101;
	mem[44] = 4'b1110;
	mem[45] = 4'b1111;
	mem[46] = 4'b1111;
	mem[47] = 4'b1111;
	mem[48] = 4'b1111;
	mem[49] = 4'b1101;
	mem[50] = 4'b1101;
	mem[51] = 4'b1110;
	mem[52] = 4'b1111;
	mem[53] = 4'b1111;
	mem[54] = 4'b1111;
	mem[55] = 4'b1111;
	mem[56] = 4'b1111;
	mem[57] = 4'b1111;
	mem[58] = 4'b1111;
	mem[59] = 4'b1111;
	mem[60] = 4'b1111;
	mem[61] = 4'b1111;
	mem[62] = 4'b1111;
	mem[63] = 4'b1111;
	mem[64] = 4'b1111;
	mem[65] = 4'b1111;
	mem[66] = 4'b1111;
	mem[67] = 4'b1111;
	mem[68] = 4'b1111;
	mem[69] = 4'b1111;
	mem[70] = 4'b1111;
	mem[71] = 4'b1001;
	mem[72] = 4'b0110;
	mem[73] = 4'b0110;
	mem[74] = 4'b0110;
	mem[75] = 4'b0110;
	mem[76] = 4'b0110;
	mem[77] = 4'b0110;
	mem[78] = 4'b0110;
	mem[79] = 4'b0110;
	mem[80] = 4'b0110;
	mem[81] = 4'b0110;
	mem[82] = 4'b0110;
	mem[83] = 4'b0111;
	mem[84] = 4'b0111;
	mem[85] = 4'b0111;
	mem[86] = 4'b0111;
	mem[87] = 4'b0111;
	mem[88] = 4'b0111;
	mem[89] = 4'b0111;
	mem[90] = 4'b0111;
	mem[91] = 4'b0111;
	mem[92] = 4'b0111;
	mem[93] = 4'b0111;
	mem[94] = 4'b0110;
	mem[95] = 4'b0110;
	mem[96] = 4'b0110;
	mem[97] = 4'b0110;
	mem[98] = 4'b0110;
	mem[99] = 4'b0111;
	mem[100] = 4'b0111;
	mem[101] = 4'b0111;
	mem[102] = 4'b0111;
	mem[103] = 4'b0111;
	mem[104] = 4'b0111;
	mem[105] = 4'b0111;
	mem[106] = 4'b0111;
	mem[107] = 4'b0111;
	mem[108] = 4'b0111;
	mem[109] = 4'b1000;
	mem[110] = 4'b0111;
	mem[111] = 4'b0111;
	mem[112] = 4'b0111;
	mem[113] = 4'b0111;
	mem[114] = 4'b0111;
	mem[115] = 4'b0111;
	mem[116] = 4'b0111;
	mem[117] = 4'b0111;
	mem[118] = 4'b0111;
	mem[119] = 4'b0111;
	mem[120] = 4'b0000;
	mem[121] = 4'b0000;
	mem[122] = 4'b0000;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b0111;
	mem[132] = 4'b1100;
	mem[133] = 4'b1101;
	mem[134] = 4'b1101;
	mem[135] = 4'b1101;
	mem[136] = 4'b1101;
	mem[137] = 4'b1101;
	mem[138] = 4'b1101;
	mem[139] = 4'b1101;
	mem[140] = 4'b1101;
	mem[141] = 4'b1101;
	mem[142] = 4'b1101;
	mem[143] = 4'b1101;
	mem[144] = 4'b1101;
	mem[145] = 4'b1101;
	mem[146] = 4'b1101;
	mem[147] = 4'b1101;
	mem[148] = 4'b1111;
	mem[149] = 4'b1111;
	mem[150] = 4'b1111;
	mem[151] = 4'b1111;
	mem[152] = 4'b1111;
	mem[153] = 4'b1111;
	mem[154] = 4'b1111;
	mem[155] = 4'b1111;
	mem[156] = 4'b1111;
	mem[157] = 4'b1111;
	mem[158] = 4'b1111;
	mem[159] = 4'b1111;
	mem[160] = 4'b1111;
	mem[161] = 4'b1111;
	mem[162] = 4'b1111;
	mem[163] = 4'b1111;
	mem[164] = 4'b1111;
	mem[165] = 4'b1111;
	mem[166] = 4'b1111;
	mem[167] = 4'b1111;
	mem[168] = 4'b1111;
	mem[169] = 4'b1111;
	mem[170] = 4'b1110;
	mem[171] = 4'b1101;
	mem[172] = 4'b1101;
	mem[173] = 4'b1110;
	mem[174] = 4'b1111;
	mem[175] = 4'b1111;
	mem[176] = 4'b1101;
	mem[177] = 4'b1101;
	mem[178] = 4'b1110;
	mem[179] = 4'b1111;
	mem[180] = 4'b1111;
	mem[181] = 4'b1111;
	mem[182] = 4'b1111;
	mem[183] = 4'b1111;
	mem[184] = 4'b1111;
	mem[185] = 4'b1111;
	mem[186] = 4'b1111;
	mem[187] = 4'b1111;
	mem[188] = 4'b1111;
	mem[189] = 4'b1111;
	mem[190] = 4'b1111;
	mem[191] = 4'b1111;
	mem[192] = 4'b1111;
	mem[193] = 4'b1111;
	mem[194] = 4'b1111;
	mem[195] = 4'b1111;
	mem[196] = 4'b1111;
	mem[197] = 4'b1111;
	mem[198] = 4'b1111;
	mem[199] = 4'b1001;
	mem[200] = 4'b0110;
	mem[201] = 4'b0110;
	mem[202] = 4'b0110;
	mem[203] = 4'b0110;
	mem[204] = 4'b0110;
	mem[205] = 4'b0110;
	mem[206] = 4'b0110;
	mem[207] = 4'b0110;
	mem[208] = 4'b0110;
	mem[209] = 4'b0110;
	mem[210] = 4'b0111;
	mem[211] = 4'b0111;
	mem[212] = 4'b0111;
	mem[213] = 4'b0111;
	mem[214] = 4'b0110;
	mem[215] = 4'b0110;
	mem[216] = 4'b0111;
	mem[217] = 4'b0111;
	mem[218] = 4'b0111;
	mem[219] = 4'b0111;
	mem[220] = 4'b0111;
	mem[221] = 4'b0111;
	mem[222] = 4'b0111;
	mem[223] = 4'b0110;
	mem[224] = 4'b0110;
	mem[225] = 4'b0110;
	mem[226] = 4'b0110;
	mem[227] = 4'b0110;
	mem[228] = 4'b0111;
	mem[229] = 4'b0111;
	mem[230] = 4'b0111;
	mem[231] = 4'b0111;
	mem[232] = 4'b0111;
	mem[233] = 4'b0111;
	mem[234] = 4'b0111;
	mem[235] = 4'b0111;
	mem[236] = 4'b1000;
	mem[237] = 4'b0111;
	mem[238] = 4'b0111;
	mem[239] = 4'b0111;
	mem[240] = 4'b0111;
	mem[241] = 4'b0111;
	mem[242] = 4'b0111;
	mem[243] = 4'b0111;
	mem[244] = 4'b0111;
	mem[245] = 4'b0111;
	mem[246] = 4'b0111;
	mem[247] = 4'b0111;
	mem[248] = 4'b0000;
	mem[249] = 4'b0000;
	mem[250] = 4'b0000;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0111;
	mem[260] = 4'b1100;
	mem[261] = 4'b1101;
	mem[262] = 4'b1101;
	mem[263] = 4'b1101;
	mem[264] = 4'b1101;
	mem[265] = 4'b1101;
	mem[266] = 4'b1101;
	mem[267] = 4'b1101;
	mem[268] = 4'b1101;
	mem[269] = 4'b1101;
	mem[270] = 4'b1101;
	mem[271] = 4'b1101;
	mem[272] = 4'b1101;
	mem[273] = 4'b1101;
	mem[274] = 4'b1101;
	mem[275] = 4'b1101;
	mem[276] = 4'b1111;
	mem[277] = 4'b1111;
	mem[278] = 4'b1111;
	mem[279] = 4'b1111;
	mem[280] = 4'b1111;
	mem[281] = 4'b1111;
	mem[282] = 4'b1111;
	mem[283] = 4'b1111;
	mem[284] = 4'b1111;
	mem[285] = 4'b1111;
	mem[286] = 4'b1111;
	mem[287] = 4'b1111;
	mem[288] = 4'b1111;
	mem[289] = 4'b1111;
	mem[290] = 4'b1111;
	mem[291] = 4'b1111;
	mem[292] = 4'b1111;
	mem[293] = 4'b1111;
	mem[294] = 4'b1111;
	mem[295] = 4'b1111;
	mem[296] = 4'b1111;
	mem[297] = 4'b1111;
	mem[298] = 4'b1111;
	mem[299] = 4'b1110;
	mem[300] = 4'b1101;
	mem[301] = 4'b1101;
	mem[302] = 4'b1110;
	mem[303] = 4'b1110;
	mem[304] = 4'b1101;
	mem[305] = 4'b1110;
	mem[306] = 4'b1111;
	mem[307] = 4'b1111;
	mem[308] = 4'b1111;
	mem[309] = 4'b1111;
	mem[310] = 4'b1111;
	mem[311] = 4'b1111;
	mem[312] = 4'b1111;
	mem[313] = 4'b1111;
	mem[314] = 4'b1111;
	mem[315] = 4'b1111;
	mem[316] = 4'b1111;
	mem[317] = 4'b1111;
	mem[318] = 4'b1111;
	mem[319] = 4'b1111;
	mem[320] = 4'b1111;
	mem[321] = 4'b1111;
	mem[322] = 4'b1111;
	mem[323] = 4'b1111;
	mem[324] = 4'b1111;
	mem[325] = 4'b1111;
	mem[326] = 4'b1111;
	mem[327] = 4'b1001;
	mem[328] = 4'b0110;
	mem[329] = 4'b0110;
	mem[330] = 4'b0110;
	mem[331] = 4'b0110;
	mem[332] = 4'b0110;
	mem[333] = 4'b0110;
	mem[334] = 4'b0110;
	mem[335] = 4'b0110;
	mem[336] = 4'b0111;
	mem[337] = 4'b0111;
	mem[338] = 4'b0111;
	mem[339] = 4'b0111;
	mem[340] = 4'b0110;
	mem[341] = 4'b0110;
	mem[342] = 4'b0110;
	mem[343] = 4'b0110;
	mem[344] = 4'b0110;
	mem[345] = 4'b0110;
	mem[346] = 4'b0111;
	mem[347] = 4'b0111;
	mem[348] = 4'b0111;
	mem[349] = 4'b0111;
	mem[350] = 4'b0111;
	mem[351] = 4'b0111;
	mem[352] = 4'b0110;
	mem[353] = 4'b0110;
	mem[354] = 4'b0110;
	mem[355] = 4'b0110;
	mem[356] = 4'b0110;
	mem[357] = 4'b0111;
	mem[358] = 4'b0111;
	mem[359] = 4'b0111;
	mem[360] = 4'b0111;
	mem[361] = 4'b0111;
	mem[362] = 4'b0111;
	mem[363] = 4'b0111;
	mem[364] = 4'b0111;
	mem[365] = 4'b0111;
	mem[366] = 4'b0111;
	mem[367] = 4'b0111;
	mem[368] = 4'b0111;
	mem[369] = 4'b0111;
	mem[370] = 4'b0111;
	mem[371] = 4'b0111;
	mem[372] = 4'b0111;
	mem[373] = 4'b0111;
	mem[374] = 4'b0111;
	mem[375] = 4'b0111;
	mem[376] = 4'b0000;
	mem[377] = 4'b0000;
	mem[378] = 4'b0000;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0111;
	mem[388] = 4'b1100;
	mem[389] = 4'b1101;
	mem[390] = 4'b1101;
	mem[391] = 4'b1101;
	mem[392] = 4'b1101;
	mem[393] = 4'b1101;
	mem[394] = 4'b1101;
	mem[395] = 4'b1101;
	mem[396] = 4'b1101;
	mem[397] = 4'b1101;
	mem[398] = 4'b1101;
	mem[399] = 4'b1101;
	mem[400] = 4'b1101;
	mem[401] = 4'b1101;
	mem[402] = 4'b1101;
	mem[403] = 4'b1101;
	mem[404] = 4'b1111;
	mem[405] = 4'b1111;
	mem[406] = 4'b1111;
	mem[407] = 4'b1111;
	mem[408] = 4'b1111;
	mem[409] = 4'b1111;
	mem[410] = 4'b1111;
	mem[411] = 4'b1111;
	mem[412] = 4'b1111;
	mem[413] = 4'b1111;
	mem[414] = 4'b1111;
	mem[415] = 4'b1111;
	mem[416] = 4'b1111;
	mem[417] = 4'b1111;
	mem[418] = 4'b1111;
	mem[419] = 4'b1111;
	mem[420] = 4'b1111;
	mem[421] = 4'b1111;
	mem[422] = 4'b1111;
	mem[423] = 4'b1111;
	mem[424] = 4'b1111;
	mem[425] = 4'b1110;
	mem[426] = 4'b1111;
	mem[427] = 4'b1111;
	mem[428] = 4'b1110;
	mem[429] = 4'b1101;
	mem[430] = 4'b1101;
	mem[431] = 4'b1101;
	mem[432] = 4'b1110;
	mem[433] = 4'b1111;
	mem[434] = 4'b1111;
	mem[435] = 4'b1111;
	mem[436] = 4'b1111;
	mem[437] = 4'b1111;
	mem[438] = 4'b1111;
	mem[439] = 4'b1111;
	mem[440] = 4'b1111;
	mem[441] = 4'b1111;
	mem[442] = 4'b1111;
	mem[443] = 4'b1111;
	mem[444] = 4'b1111;
	mem[445] = 4'b1111;
	mem[446] = 4'b1111;
	mem[447] = 4'b1111;
	mem[448] = 4'b1111;
	mem[449] = 4'b1111;
	mem[450] = 4'b1111;
	mem[451] = 4'b1111;
	mem[452] = 4'b1111;
	mem[453] = 4'b1111;
	mem[454] = 4'b1111;
	mem[455] = 4'b1001;
	mem[456] = 4'b0110;
	mem[457] = 4'b0110;
	mem[458] = 4'b0110;
	mem[459] = 4'b0110;
	mem[460] = 4'b0110;
	mem[461] = 4'b0110;
	mem[462] = 4'b0111;
	mem[463] = 4'b0111;
	mem[464] = 4'b0111;
	mem[465] = 4'b0111;
	mem[466] = 4'b0111;
	mem[467] = 4'b0110;
	mem[468] = 4'b0110;
	mem[469] = 4'b0110;
	mem[470] = 4'b0110;
	mem[471] = 4'b0110;
	mem[472] = 4'b0110;
	mem[473] = 4'b0110;
	mem[474] = 4'b0110;
	mem[475] = 4'b0111;
	mem[476] = 4'b0111;
	mem[477] = 4'b0111;
	mem[478] = 4'b0111;
	mem[479] = 4'b0111;
	mem[480] = 4'b0111;
	mem[481] = 4'b0110;
	mem[482] = 4'b0110;
	mem[483] = 4'b0110;
	mem[484] = 4'b0110;
	mem[485] = 4'b0110;
	mem[486] = 4'b0111;
	mem[487] = 4'b0111;
	mem[488] = 4'b0111;
	mem[489] = 4'b0111;
	mem[490] = 4'b0111;
	mem[491] = 4'b0111;
	mem[492] = 4'b0111;
	mem[493] = 4'b0111;
	mem[494] = 4'b0111;
	mem[495] = 4'b0111;
	mem[496] = 4'b0111;
	mem[497] = 4'b0111;
	mem[498] = 4'b0111;
	mem[499] = 4'b0111;
	mem[500] = 4'b0111;
	mem[501] = 4'b0111;
	mem[502] = 4'b0111;
	mem[503] = 4'b0111;
	mem[504] = 4'b0000;
	mem[505] = 4'b0000;
	mem[506] = 4'b0000;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0111;
	mem[516] = 4'b1100;
	mem[517] = 4'b1101;
	mem[518] = 4'b1101;
	mem[519] = 4'b1101;
	mem[520] = 4'b1101;
	mem[521] = 4'b1101;
	mem[522] = 4'b1101;
	mem[523] = 4'b1101;
	mem[524] = 4'b1101;
	mem[525] = 4'b1101;
	mem[526] = 4'b1101;
	mem[527] = 4'b1101;
	mem[528] = 4'b1101;
	mem[529] = 4'b1101;
	mem[530] = 4'b1101;
	mem[531] = 4'b1101;
	mem[532] = 4'b1111;
	mem[533] = 4'b1111;
	mem[534] = 4'b1111;
	mem[535] = 4'b1111;
	mem[536] = 4'b1111;
	mem[537] = 4'b1111;
	mem[538] = 4'b1111;
	mem[539] = 4'b1111;
	mem[540] = 4'b1111;
	mem[541] = 4'b1111;
	mem[542] = 4'b1111;
	mem[543] = 4'b1111;
	mem[544] = 4'b1111;
	mem[545] = 4'b1111;
	mem[546] = 4'b1111;
	mem[547] = 4'b1111;
	mem[548] = 4'b1111;
	mem[549] = 4'b1111;
	mem[550] = 4'b1111;
	mem[551] = 4'b1111;
	mem[552] = 4'b1101;
	mem[553] = 4'b1101;
	mem[554] = 4'b1110;
	mem[555] = 4'b1111;
	mem[556] = 4'b1111;
	mem[557] = 4'b1110;
	mem[558] = 4'b1101;
	mem[559] = 4'b1110;
	mem[560] = 4'b1111;
	mem[561] = 4'b1111;
	mem[562] = 4'b1111;
	mem[563] = 4'b1111;
	mem[564] = 4'b1111;
	mem[565] = 4'b1111;
	mem[566] = 4'b1111;
	mem[567] = 4'b1111;
	mem[568] = 4'b1111;
	mem[569] = 4'b1111;
	mem[570] = 4'b1111;
	mem[571] = 4'b1111;
	mem[572] = 4'b1111;
	mem[573] = 4'b1111;
	mem[574] = 4'b1111;
	mem[575] = 4'b1111;
	mem[576] = 4'b1111;
	mem[577] = 4'b1111;
	mem[578] = 4'b1111;
	mem[579] = 4'b1111;
	mem[580] = 4'b1111;
	mem[581] = 4'b1111;
	mem[582] = 4'b1111;
	mem[583] = 4'b1001;
	mem[584] = 4'b0110;
	mem[585] = 4'b0110;
	mem[586] = 4'b0110;
	mem[587] = 4'b0110;
	mem[588] = 4'b0111;
	mem[589] = 4'b0111;
	mem[590] = 4'b0111;
	mem[591] = 4'b0111;
	mem[592] = 4'b0111;
	mem[593] = 4'b0111;
	mem[594] = 4'b0110;
	mem[595] = 4'b0110;
	mem[596] = 4'b0110;
	mem[597] = 4'b0110;
	mem[598] = 4'b0110;
	mem[599] = 4'b0110;
	mem[600] = 4'b0110;
	mem[601] = 4'b0110;
	mem[602] = 4'b0110;
	mem[603] = 4'b0110;
	mem[604] = 4'b0111;
	mem[605] = 4'b0111;
	mem[606] = 4'b0111;
	mem[607] = 4'b0111;
	mem[608] = 4'b0111;
	mem[609] = 4'b0111;
	mem[610] = 4'b0110;
	mem[611] = 4'b0110;
	mem[612] = 4'b0110;
	mem[613] = 4'b0110;
	mem[614] = 4'b0111;
	mem[615] = 4'b0111;
	mem[616] = 4'b0111;
	mem[617] = 4'b0111;
	mem[618] = 4'b0111;
	mem[619] = 4'b0111;
	mem[620] = 4'b0111;
	mem[621] = 4'b0111;
	mem[622] = 4'b0111;
	mem[623] = 4'b0111;
	mem[624] = 4'b0111;
	mem[625] = 4'b0111;
	mem[626] = 4'b0111;
	mem[627] = 4'b0111;
	mem[628] = 4'b0111;
	mem[629] = 4'b0111;
	mem[630] = 4'b0111;
	mem[631] = 4'b0111;
	mem[632] = 4'b0000;
	mem[633] = 4'b0000;
	mem[634] = 4'b0000;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0111;
	mem[644] = 4'b1100;
	mem[645] = 4'b1101;
	mem[646] = 4'b1101;
	mem[647] = 4'b1101;
	mem[648] = 4'b1101;
	mem[649] = 4'b1101;
	mem[650] = 4'b1101;
	mem[651] = 4'b1101;
	mem[652] = 4'b1101;
	mem[653] = 4'b1101;
	mem[654] = 4'b1101;
	mem[655] = 4'b1101;
	mem[656] = 4'b1101;
	mem[657] = 4'b1101;
	mem[658] = 4'b1101;
	mem[659] = 4'b1101;
	mem[660] = 4'b1111;
	mem[661] = 4'b1111;
	mem[662] = 4'b1111;
	mem[663] = 4'b1111;
	mem[664] = 4'b1111;
	mem[665] = 4'b1111;
	mem[666] = 4'b1111;
	mem[667] = 4'b1111;
	mem[668] = 4'b1111;
	mem[669] = 4'b1111;
	mem[670] = 4'b1111;
	mem[671] = 4'b1111;
	mem[672] = 4'b1111;
	mem[673] = 4'b1111;
	mem[674] = 4'b1111;
	mem[675] = 4'b1111;
	mem[676] = 4'b1111;
	mem[677] = 4'b1111;
	mem[678] = 4'b1111;
	mem[679] = 4'b1101;
	mem[680] = 4'b1101;
	mem[681] = 4'b1110;
	mem[682] = 4'b1111;
	mem[683] = 4'b1111;
	mem[684] = 4'b1111;
	mem[685] = 4'b1111;
	mem[686] = 4'b1111;
	mem[687] = 4'b1111;
	mem[688] = 4'b1111;
	mem[689] = 4'b1111;
	mem[690] = 4'b1111;
	mem[691] = 4'b1111;
	mem[692] = 4'b1111;
	mem[693] = 4'b1111;
	mem[694] = 4'b1111;
	mem[695] = 4'b1111;
	mem[696] = 4'b1111;
	mem[697] = 4'b1111;
	mem[698] = 4'b1111;
	mem[699] = 4'b1111;
	mem[700] = 4'b1111;
	mem[701] = 4'b1111;
	mem[702] = 4'b1111;
	mem[703] = 4'b1111;
	mem[704] = 4'b1111;
	mem[705] = 4'b1111;
	mem[706] = 4'b1111;
	mem[707] = 4'b1111;
	mem[708] = 4'b1111;
	mem[709] = 4'b1111;
	mem[710] = 4'b1111;
	mem[711] = 4'b1001;
	mem[712] = 4'b0110;
	mem[713] = 4'b0110;
	mem[714] = 4'b0111;
	mem[715] = 4'b0111;
	mem[716] = 4'b0111;
	mem[717] = 4'b0111;
	mem[718] = 4'b0111;
	mem[719] = 4'b0111;
	mem[720] = 4'b0111;
	mem[721] = 4'b0110;
	mem[722] = 4'b0110;
	mem[723] = 4'b0110;
	mem[724] = 4'b0110;
	mem[725] = 4'b0111;
	mem[726] = 4'b0111;
	mem[727] = 4'b0111;
	mem[728] = 4'b0110;
	mem[729] = 4'b0110;
	mem[730] = 4'b0110;
	mem[731] = 4'b0110;
	mem[732] = 4'b0110;
	mem[733] = 4'b0111;
	mem[734] = 4'b0111;
	mem[735] = 4'b0111;
	mem[736] = 4'b0111;
	mem[737] = 4'b0111;
	mem[738] = 4'b0111;
	mem[739] = 4'b0110;
	mem[740] = 4'b0110;
	mem[741] = 4'b0110;
	mem[742] = 4'b0110;
	mem[743] = 4'b0111;
	mem[744] = 4'b0111;
	mem[745] = 4'b0111;
	mem[746] = 4'b0111;
	mem[747] = 4'b0111;
	mem[748] = 4'b0111;
	mem[749] = 4'b0111;
	mem[750] = 4'b0111;
	mem[751] = 4'b0111;
	mem[752] = 4'b0111;
	mem[753] = 4'b0111;
	mem[754] = 4'b0111;
	mem[755] = 4'b0111;
	mem[756] = 4'b0111;
	mem[757] = 4'b0111;
	mem[758] = 4'b1000;
	mem[759] = 4'b1000;
	mem[760] = 4'b0000;
	mem[761] = 4'b0000;
	mem[762] = 4'b0000;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0111;
	mem[772] = 4'b1100;
	mem[773] = 4'b1101;
	mem[774] = 4'b1101;
	mem[775] = 4'b1101;
	mem[776] = 4'b1101;
	mem[777] = 4'b1101;
	mem[778] = 4'b1101;
	mem[779] = 4'b1101;
	mem[780] = 4'b1101;
	mem[781] = 4'b1101;
	mem[782] = 4'b1101;
	mem[783] = 4'b1101;
	mem[784] = 4'b1101;
	mem[785] = 4'b1101;
	mem[786] = 4'b1101;
	mem[787] = 4'b1101;
	mem[788] = 4'b1111;
	mem[789] = 4'b1111;
	mem[790] = 4'b1111;
	mem[791] = 4'b1111;
	mem[792] = 4'b1111;
	mem[793] = 4'b1111;
	mem[794] = 4'b1111;
	mem[795] = 4'b1111;
	mem[796] = 4'b1111;
	mem[797] = 4'b1111;
	mem[798] = 4'b1111;
	mem[799] = 4'b1111;
	mem[800] = 4'b1111;
	mem[801] = 4'b1110;
	mem[802] = 4'b1110;
	mem[803] = 4'b1110;
	mem[804] = 4'b1111;
	mem[805] = 4'b1111;
	mem[806] = 4'b1111;
	mem[807] = 4'b1101;
	mem[808] = 4'b1110;
	mem[809] = 4'b1111;
	mem[810] = 4'b1111;
	mem[811] = 4'b1111;
	mem[812] = 4'b1111;
	mem[813] = 4'b1111;
	mem[814] = 4'b1111;
	mem[815] = 4'b1111;
	mem[816] = 4'b1111;
	mem[817] = 4'b1111;
	mem[818] = 4'b1111;
	mem[819] = 4'b1111;
	mem[820] = 4'b1111;
	mem[821] = 4'b1111;
	mem[822] = 4'b1111;
	mem[823] = 4'b1111;
	mem[824] = 4'b1111;
	mem[825] = 4'b1111;
	mem[826] = 4'b1111;
	mem[827] = 4'b1111;
	mem[828] = 4'b1111;
	mem[829] = 4'b1111;
	mem[830] = 4'b1111;
	mem[831] = 4'b1111;
	mem[832] = 4'b1111;
	mem[833] = 4'b1111;
	mem[834] = 4'b1111;
	mem[835] = 4'b1111;
	mem[836] = 4'b1111;
	mem[837] = 4'b1111;
	mem[838] = 4'b1111;
	mem[839] = 4'b1001;
	mem[840] = 4'b0111;
	mem[841] = 4'b0111;
	mem[842] = 4'b0111;
	mem[843] = 4'b0111;
	mem[844] = 4'b0111;
	mem[845] = 4'b0111;
	mem[846] = 4'b0111;
	mem[847] = 4'b0111;
	mem[848] = 4'b0111;
	mem[849] = 4'b0110;
	mem[850] = 4'b0110;
	mem[851] = 4'b0110;
	mem[852] = 4'b0111;
	mem[853] = 4'b1000;
	mem[854] = 4'b0111;
	mem[855] = 4'b0111;
	mem[856] = 4'b0111;
	mem[857] = 4'b0110;
	mem[858] = 4'b0110;
	mem[859] = 4'b0110;
	mem[860] = 4'b0110;
	mem[861] = 4'b0110;
	mem[862] = 4'b0111;
	mem[863] = 4'b0111;
	mem[864] = 4'b0111;
	mem[865] = 4'b0111;
	mem[866] = 4'b0111;
	mem[867] = 4'b0111;
	mem[868] = 4'b0110;
	mem[869] = 4'b0110;
	mem[870] = 4'b0111;
	mem[871] = 4'b1000;
	mem[872] = 4'b0111;
	mem[873] = 4'b0111;
	mem[874] = 4'b0111;
	mem[875] = 4'b0111;
	mem[876] = 4'b0111;
	mem[877] = 4'b0111;
	mem[878] = 4'b0110;
	mem[879] = 4'b0101;
	mem[880] = 4'b0100;
	mem[881] = 4'b0100;
	mem[882] = 4'b0011;
	mem[883] = 4'b0010;
	mem[884] = 4'b0010;
	mem[885] = 4'b0001;
	mem[886] = 4'b0000;
	mem[887] = 4'b0000;
	mem[888] = 4'b0000;
	mem[889] = 4'b0000;
	mem[890] = 4'b0000;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0111;
	mem[900] = 4'b1100;
	mem[901] = 4'b1101;
	mem[902] = 4'b1101;
	mem[903] = 4'b1101;
	mem[904] = 4'b1101;
	mem[905] = 4'b1101;
	mem[906] = 4'b1101;
	mem[907] = 4'b1101;
	mem[908] = 4'b1101;
	mem[909] = 4'b1101;
	mem[910] = 4'b1101;
	mem[911] = 4'b1101;
	mem[912] = 4'b1101;
	mem[913] = 4'b1101;
	mem[914] = 4'b1101;
	mem[915] = 4'b1101;
	mem[916] = 4'b1111;
	mem[917] = 4'b1111;
	mem[918] = 4'b1111;
	mem[919] = 4'b1111;
	mem[920] = 4'b1111;
	mem[921] = 4'b1111;
	mem[922] = 4'b1111;
	mem[923] = 4'b1111;
	mem[924] = 4'b1111;
	mem[925] = 4'b1111;
	mem[926] = 4'b1111;
	mem[927] = 4'b1111;
	mem[928] = 4'b1110;
	mem[929] = 4'b1101;
	mem[930] = 4'b1101;
	mem[931] = 4'b1111;
	mem[932] = 4'b1111;
	mem[933] = 4'b1111;
	mem[934] = 4'b1111;
	mem[935] = 4'b1111;
	mem[936] = 4'b1111;
	mem[937] = 4'b1111;
	mem[938] = 4'b1111;
	mem[939] = 4'b1111;
	mem[940] = 4'b1111;
	mem[941] = 4'b1111;
	mem[942] = 4'b1111;
	mem[943] = 4'b1111;
	mem[944] = 4'b1111;
	mem[945] = 4'b1111;
	mem[946] = 4'b1111;
	mem[947] = 4'b1111;
	mem[948] = 4'b1111;
	mem[949] = 4'b1111;
	mem[950] = 4'b1111;
	mem[951] = 4'b1111;
	mem[952] = 4'b1111;
	mem[953] = 4'b1111;
	mem[954] = 4'b1111;
	mem[955] = 4'b1111;
	mem[956] = 4'b1111;
	mem[957] = 4'b1111;
	mem[958] = 4'b1111;
	mem[959] = 4'b1111;
	mem[960] = 4'b1111;
	mem[961] = 4'b1111;
	mem[962] = 4'b1111;
	mem[963] = 4'b1111;
	mem[964] = 4'b1111;
	mem[965] = 4'b1111;
	mem[966] = 4'b1111;
	mem[967] = 4'b1001;
	mem[968] = 4'b0111;
	mem[969] = 4'b0111;
	mem[970] = 4'b0111;
	mem[971] = 4'b0111;
	mem[972] = 4'b0111;
	mem[973] = 4'b0111;
	mem[974] = 4'b0111;
	mem[975] = 4'b0111;
	mem[976] = 4'b0110;
	mem[977] = 4'b0110;
	mem[978] = 4'b0110;
	mem[979] = 4'b0110;
	mem[980] = 4'b1000;
	mem[981] = 4'b0111;
	mem[982] = 4'b0111;
	mem[983] = 4'b0111;
	mem[984] = 4'b0110;
	mem[985] = 4'b0110;
	mem[986] = 4'b0110;
	mem[987] = 4'b0110;
	mem[988] = 4'b0110;
	mem[989] = 4'b0110;
	mem[990] = 4'b0110;
	mem[991] = 4'b0111;
	mem[992] = 4'b0111;
	mem[993] = 4'b0111;
	mem[994] = 4'b0111;
	mem[995] = 4'b0111;
	mem[996] = 4'b0111;
	mem[997] = 4'b0111;
	mem[998] = 4'b0111;
	mem[999] = 4'b0101;
	mem[1000] = 4'b0100;
	mem[1001] = 4'b0011;
	mem[1002] = 4'b0010;
	mem[1003] = 4'b0001;
	mem[1004] = 4'b0000;
	mem[1005] = 4'b0000;
	mem[1006] = 4'b0000;
	mem[1007] = 4'b0000;
	mem[1008] = 4'b0000;
	mem[1009] = 4'b0000;
	mem[1010] = 4'b0000;
	mem[1011] = 4'b0000;
	mem[1012] = 4'b0000;
	mem[1013] = 4'b0000;
	mem[1014] = 4'b0000;
	mem[1015] = 4'b0000;
	mem[1016] = 4'b0000;
	mem[1017] = 4'b0000;
	mem[1018] = 4'b0000;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0111;
	mem[1028] = 4'b1100;
	mem[1029] = 4'b1101;
	mem[1030] = 4'b1101;
	mem[1031] = 4'b1101;
	mem[1032] = 4'b1101;
	mem[1033] = 4'b1101;
	mem[1034] = 4'b1101;
	mem[1035] = 4'b1101;
	mem[1036] = 4'b1101;
	mem[1037] = 4'b1101;
	mem[1038] = 4'b1101;
	mem[1039] = 4'b1101;
	mem[1040] = 4'b1101;
	mem[1041] = 4'b1101;
	mem[1042] = 4'b1101;
	mem[1043] = 4'b1101;
	mem[1044] = 4'b1111;
	mem[1045] = 4'b1111;
	mem[1046] = 4'b1111;
	mem[1047] = 4'b1111;
	mem[1048] = 4'b1111;
	mem[1049] = 4'b1111;
	mem[1050] = 4'b1111;
	mem[1051] = 4'b1111;
	mem[1052] = 4'b1111;
	mem[1053] = 4'b1111;
	mem[1054] = 4'b1111;
	mem[1055] = 4'b1110;
	mem[1056] = 4'b1101;
	mem[1057] = 4'b1111;
	mem[1058] = 4'b1111;
	mem[1059] = 4'b1111;
	mem[1060] = 4'b1111;
	mem[1061] = 4'b1110;
	mem[1062] = 4'b1111;
	mem[1063] = 4'b1111;
	mem[1064] = 4'b1111;
	mem[1065] = 4'b1111;
	mem[1066] = 4'b1111;
	mem[1067] = 4'b1111;
	mem[1068] = 4'b1111;
	mem[1069] = 4'b1111;
	mem[1070] = 4'b1111;
	mem[1071] = 4'b1111;
	mem[1072] = 4'b1111;
	mem[1073] = 4'b1111;
	mem[1074] = 4'b1111;
	mem[1075] = 4'b1111;
	mem[1076] = 4'b1111;
	mem[1077] = 4'b1111;
	mem[1078] = 4'b1111;
	mem[1079] = 4'b1111;
	mem[1080] = 4'b1111;
	mem[1081] = 4'b1111;
	mem[1082] = 4'b1111;
	mem[1083] = 4'b1111;
	mem[1084] = 4'b1111;
	mem[1085] = 4'b1111;
	mem[1086] = 4'b1111;
	mem[1087] = 4'b1111;
	mem[1088] = 4'b1111;
	mem[1089] = 4'b1111;
	mem[1090] = 4'b1111;
	mem[1091] = 4'b1111;
	mem[1092] = 4'b1111;
	mem[1093] = 4'b1111;
	mem[1094] = 4'b1111;
	mem[1095] = 4'b1001;
	mem[1096] = 4'b0111;
	mem[1097] = 4'b0111;
	mem[1098] = 4'b0111;
	mem[1099] = 4'b0111;
	mem[1100] = 4'b0111;
	mem[1101] = 4'b0111;
	mem[1102] = 4'b0111;
	mem[1103] = 4'b0111;
	mem[1104] = 4'b0110;
	mem[1105] = 4'b0110;
	mem[1106] = 4'b0110;
	mem[1107] = 4'b0111;
	mem[1108] = 4'b0111;
	mem[1109] = 4'b0111;
	mem[1110] = 4'b0111;
	mem[1111] = 4'b0110;
	mem[1112] = 4'b0110;
	mem[1113] = 4'b0111;
	mem[1114] = 4'b0111;
	mem[1115] = 4'b0110;
	mem[1116] = 4'b0110;
	mem[1117] = 4'b0110;
	mem[1118] = 4'b0110;
	mem[1119] = 4'b0110;
	mem[1120] = 4'b0110;
	mem[1121] = 4'b0101;
	mem[1122] = 4'b0011;
	mem[1123] = 4'b0010;
	mem[1124] = 4'b0001;
	mem[1125] = 4'b0001;
	mem[1126] = 4'b0000;
	mem[1127] = 4'b0000;
	mem[1128] = 4'b0000;
	mem[1129] = 4'b0000;
	mem[1130] = 4'b0000;
	mem[1131] = 4'b0000;
	mem[1132] = 4'b0000;
	mem[1133] = 4'b0000;
	mem[1134] = 4'b0000;
	mem[1135] = 4'b0000;
	mem[1136] = 4'b0000;
	mem[1137] = 4'b0000;
	mem[1138] = 4'b0000;
	mem[1139] = 4'b0000;
	mem[1140] = 4'b0000;
	mem[1141] = 4'b0000;
	mem[1142] = 4'b0000;
	mem[1143] = 4'b0000;
	mem[1144] = 4'b0000;
	mem[1145] = 4'b0000;
	mem[1146] = 4'b0000;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0111;
	mem[1156] = 4'b1100;
	mem[1157] = 4'b1101;
	mem[1158] = 4'b1101;
	mem[1159] = 4'b1101;
	mem[1160] = 4'b1101;
	mem[1161] = 4'b1101;
	mem[1162] = 4'b1101;
	mem[1163] = 4'b1101;
	mem[1164] = 4'b1101;
	mem[1165] = 4'b1101;
	mem[1166] = 4'b1101;
	mem[1167] = 4'b1101;
	mem[1168] = 4'b1101;
	mem[1169] = 4'b1101;
	mem[1170] = 4'b1101;
	mem[1171] = 4'b1101;
	mem[1172] = 4'b1111;
	mem[1173] = 4'b1111;
	mem[1174] = 4'b1111;
	mem[1175] = 4'b1111;
	mem[1176] = 4'b1111;
	mem[1177] = 4'b1111;
	mem[1178] = 4'b1111;
	mem[1179] = 4'b1111;
	mem[1180] = 4'b1111;
	mem[1181] = 4'b1111;
	mem[1182] = 4'b1110;
	mem[1183] = 4'b1101;
	mem[1184] = 4'b1111;
	mem[1185] = 4'b1111;
	mem[1186] = 4'b1111;
	mem[1187] = 4'b1110;
	mem[1188] = 4'b1101;
	mem[1189] = 4'b1101;
	mem[1190] = 4'b1101;
	mem[1191] = 4'b1111;
	mem[1192] = 4'b1111;
	mem[1193] = 4'b1111;
	mem[1194] = 4'b1111;
	mem[1195] = 4'b1111;
	mem[1196] = 4'b1111;
	mem[1197] = 4'b1111;
	mem[1198] = 4'b1111;
	mem[1199] = 4'b1111;
	mem[1200] = 4'b1111;
	mem[1201] = 4'b1111;
	mem[1202] = 4'b1111;
	mem[1203] = 4'b1111;
	mem[1204] = 4'b1111;
	mem[1205] = 4'b1111;
	mem[1206] = 4'b1111;
	mem[1207] = 4'b1111;
	mem[1208] = 4'b1111;
	mem[1209] = 4'b1111;
	mem[1210] = 4'b1111;
	mem[1211] = 4'b1111;
	mem[1212] = 4'b1111;
	mem[1213] = 4'b1111;
	mem[1214] = 4'b1111;
	mem[1215] = 4'b1111;
	mem[1216] = 4'b1111;
	mem[1217] = 4'b1111;
	mem[1218] = 4'b1111;
	mem[1219] = 4'b1111;
	mem[1220] = 4'b1111;
	mem[1221] = 4'b1111;
	mem[1222] = 4'b1111;
	mem[1223] = 4'b1001;
	mem[1224] = 4'b0111;
	mem[1225] = 4'b0111;
	mem[1226] = 4'b0111;
	mem[1227] = 4'b0111;
	mem[1228] = 4'b0111;
	mem[1229] = 4'b0111;
	mem[1230] = 4'b0111;
	mem[1231] = 4'b0111;
	mem[1232] = 4'b0111;
	mem[1233] = 4'b0110;
	mem[1234] = 4'b0110;
	mem[1235] = 4'b0111;
	mem[1236] = 4'b1000;
	mem[1237] = 4'b0111;
	mem[1238] = 4'b0111;
	mem[1239] = 4'b0110;
	mem[1240] = 4'b0110;
	mem[1241] = 4'b1000;
	mem[1242] = 4'b0111;
	mem[1243] = 4'b0101;
	mem[1244] = 4'b0011;
	mem[1245] = 4'b0010;
	mem[1246] = 4'b0001;
	mem[1247] = 4'b0000;
	mem[1248] = 4'b0000;
	mem[1249] = 4'b0000;
	mem[1250] = 4'b0000;
	mem[1251] = 4'b0000;
	mem[1252] = 4'b0000;
	mem[1253] = 4'b0000;
	mem[1254] = 4'b0000;
	mem[1255] = 4'b0000;
	mem[1256] = 4'b0000;
	mem[1257] = 4'b0000;
	mem[1258] = 4'b0000;
	mem[1259] = 4'b0000;
	mem[1260] = 4'b0000;
	mem[1261] = 4'b0000;
	mem[1262] = 4'b0000;
	mem[1263] = 4'b0000;
	mem[1264] = 4'b0000;
	mem[1265] = 4'b0000;
	mem[1266] = 4'b0000;
	mem[1267] = 4'b0000;
	mem[1268] = 4'b0000;
	mem[1269] = 4'b0000;
	mem[1270] = 4'b0000;
	mem[1271] = 4'b0000;
	mem[1272] = 4'b0000;
	mem[1273] = 4'b0000;
	mem[1274] = 4'b0000;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0111;
	mem[1284] = 4'b1100;
	mem[1285] = 4'b1101;
	mem[1286] = 4'b1101;
	mem[1287] = 4'b1101;
	mem[1288] = 4'b1101;
	mem[1289] = 4'b1101;
	mem[1290] = 4'b1101;
	mem[1291] = 4'b1101;
	mem[1292] = 4'b1101;
	mem[1293] = 4'b1101;
	mem[1294] = 4'b1101;
	mem[1295] = 4'b1101;
	mem[1296] = 4'b1101;
	mem[1297] = 4'b1101;
	mem[1298] = 4'b1101;
	mem[1299] = 4'b1101;
	mem[1300] = 4'b1111;
	mem[1301] = 4'b1111;
	mem[1302] = 4'b1111;
	mem[1303] = 4'b1111;
	mem[1304] = 4'b1111;
	mem[1305] = 4'b1111;
	mem[1306] = 4'b1111;
	mem[1307] = 4'b1111;
	mem[1308] = 4'b1111;
	mem[1309] = 4'b1111;
	mem[1310] = 4'b1110;
	mem[1311] = 4'b1101;
	mem[1312] = 4'b1110;
	mem[1313] = 4'b1110;
	mem[1314] = 4'b1101;
	mem[1315] = 4'b1101;
	mem[1316] = 4'b1110;
	mem[1317] = 4'b1110;
	mem[1318] = 4'b1101;
	mem[1319] = 4'b1110;
	mem[1320] = 4'b1111;
	mem[1321] = 4'b1111;
	mem[1322] = 4'b1111;
	mem[1323] = 4'b1111;
	mem[1324] = 4'b1111;
	mem[1325] = 4'b1111;
	mem[1326] = 4'b1111;
	mem[1327] = 4'b1111;
	mem[1328] = 4'b1111;
	mem[1329] = 4'b1111;
	mem[1330] = 4'b1111;
	mem[1331] = 4'b1111;
	mem[1332] = 4'b1111;
	mem[1333] = 4'b1111;
	mem[1334] = 4'b1111;
	mem[1335] = 4'b1111;
	mem[1336] = 4'b1111;
	mem[1337] = 4'b1111;
	mem[1338] = 4'b1111;
	mem[1339] = 4'b1111;
	mem[1340] = 4'b1111;
	mem[1341] = 4'b1111;
	mem[1342] = 4'b1111;
	mem[1343] = 4'b1111;
	mem[1344] = 4'b1111;
	mem[1345] = 4'b1111;
	mem[1346] = 4'b1111;
	mem[1347] = 4'b1111;
	mem[1348] = 4'b1111;
	mem[1349] = 4'b1111;
	mem[1350] = 4'b1111;
	mem[1351] = 4'b1001;
	mem[1352] = 4'b0111;
	mem[1353] = 4'b0111;
	mem[1354] = 4'b0111;
	mem[1355] = 4'b0111;
	mem[1356] = 4'b0111;
	mem[1357] = 4'b0111;
	mem[1358] = 4'b0111;
	mem[1359] = 4'b0111;
	mem[1360] = 4'b0111;
	mem[1361] = 4'b0110;
	mem[1362] = 4'b0111;
	mem[1363] = 4'b1000;
	mem[1364] = 4'b0111;
	mem[1365] = 4'b0110;
	mem[1366] = 4'b0100;
	mem[1367] = 4'b0011;
	mem[1368] = 4'b0010;
	mem[1369] = 4'b0001;
	mem[1370] = 4'b0000;
	mem[1371] = 4'b0000;
	mem[1372] = 4'b0000;
	mem[1373] = 4'b0000;
	mem[1374] = 4'b0000;
	mem[1375] = 4'b0000;
	mem[1376] = 4'b0000;
	mem[1377] = 4'b0000;
	mem[1378] = 4'b0001;
	mem[1379] = 4'b0000;
	mem[1380] = 4'b0000;
	mem[1381] = 4'b0000;
	mem[1382] = 4'b0000;
	mem[1383] = 4'b0000;
	mem[1384] = 4'b0000;
	mem[1385] = 4'b0000;
	mem[1386] = 4'b0000;
	mem[1387] = 4'b0000;
	mem[1388] = 4'b0000;
	mem[1389] = 4'b0000;
	mem[1390] = 4'b0000;
	mem[1391] = 4'b0000;
	mem[1392] = 4'b0000;
	mem[1393] = 4'b0000;
	mem[1394] = 4'b0000;
	mem[1395] = 4'b0000;
	mem[1396] = 4'b0000;
	mem[1397] = 4'b0000;
	mem[1398] = 4'b0000;
	mem[1399] = 4'b0000;
	mem[1400] = 4'b0000;
	mem[1401] = 4'b0000;
	mem[1402] = 4'b0000;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0111;
	mem[1412] = 4'b1100;
	mem[1413] = 4'b1101;
	mem[1414] = 4'b1101;
	mem[1415] = 4'b1101;
	mem[1416] = 4'b1101;
	mem[1417] = 4'b1101;
	mem[1418] = 4'b1101;
	mem[1419] = 4'b1101;
	mem[1420] = 4'b1101;
	mem[1421] = 4'b1101;
	mem[1422] = 4'b1101;
	mem[1423] = 4'b1101;
	mem[1424] = 4'b1101;
	mem[1425] = 4'b1101;
	mem[1426] = 4'b1101;
	mem[1427] = 4'b1101;
	mem[1428] = 4'b1111;
	mem[1429] = 4'b1111;
	mem[1430] = 4'b1111;
	mem[1431] = 4'b1111;
	mem[1432] = 4'b1111;
	mem[1433] = 4'b1111;
	mem[1434] = 4'b1111;
	mem[1435] = 4'b1111;
	mem[1436] = 4'b1111;
	mem[1437] = 4'b1111;
	mem[1438] = 4'b1111;
	mem[1439] = 4'b1101;
	mem[1440] = 4'b1101;
	mem[1441] = 4'b1101;
	mem[1442] = 4'b1101;
	mem[1443] = 4'b1110;
	mem[1444] = 4'b1111;
	mem[1445] = 4'b1111;
	mem[1446] = 4'b1101;
	mem[1447] = 4'b1110;
	mem[1448] = 4'b1111;
	mem[1449] = 4'b1111;
	mem[1450] = 4'b1111;
	mem[1451] = 4'b1111;
	mem[1452] = 4'b1111;
	mem[1453] = 4'b1111;
	mem[1454] = 4'b1111;
	mem[1455] = 4'b1111;
	mem[1456] = 4'b1111;
	mem[1457] = 4'b1111;
	mem[1458] = 4'b1111;
	mem[1459] = 4'b1111;
	mem[1460] = 4'b1111;
	mem[1461] = 4'b1111;
	mem[1462] = 4'b1111;
	mem[1463] = 4'b1111;
	mem[1464] = 4'b1111;
	mem[1465] = 4'b1111;
	mem[1466] = 4'b1111;
	mem[1467] = 4'b1111;
	mem[1468] = 4'b1111;
	mem[1469] = 4'b1111;
	mem[1470] = 4'b1111;
	mem[1471] = 4'b1111;
	mem[1472] = 4'b1111;
	mem[1473] = 4'b1111;
	mem[1474] = 4'b1111;
	mem[1475] = 4'b1111;
	mem[1476] = 4'b1111;
	mem[1477] = 4'b1111;
	mem[1478] = 4'b1111;
	mem[1479] = 4'b1001;
	mem[1480] = 4'b0111;
	mem[1481] = 4'b0111;
	mem[1482] = 4'b0111;
	mem[1483] = 4'b0111;
	mem[1484] = 4'b0111;
	mem[1485] = 4'b0111;
	mem[1486] = 4'b0111;
	mem[1487] = 4'b0111;
	mem[1488] = 4'b0111;
	mem[1489] = 4'b0110;
	mem[1490] = 4'b0100;
	mem[1491] = 4'b0010;
	mem[1492] = 4'b0000;
	mem[1493] = 4'b0000;
	mem[1494] = 4'b0000;
	mem[1495] = 4'b0000;
	mem[1496] = 4'b0001;
	mem[1497] = 4'b0000;
	mem[1498] = 4'b0000;
	mem[1499] = 4'b0000;
	mem[1500] = 4'b0000;
	mem[1501] = 4'b0000;
	mem[1502] = 4'b0000;
	mem[1503] = 4'b0000;
	mem[1504] = 4'b0000;
	mem[1505] = 4'b0001;
	mem[1506] = 4'b0000;
	mem[1507] = 4'b0000;
	mem[1508] = 4'b0000;
	mem[1509] = 4'b0000;
	mem[1510] = 4'b0000;
	mem[1511] = 4'b0000;
	mem[1512] = 4'b0000;
	mem[1513] = 4'b0000;
	mem[1514] = 4'b0000;
	mem[1515] = 4'b0000;
	mem[1516] = 4'b0000;
	mem[1517] = 4'b0000;
	mem[1518] = 4'b0000;
	mem[1519] = 4'b0000;
	mem[1520] = 4'b0000;
	mem[1521] = 4'b0000;
	mem[1522] = 4'b0000;
	mem[1523] = 4'b0000;
	mem[1524] = 4'b0000;
	mem[1525] = 4'b0000;
	mem[1526] = 4'b0000;
	mem[1527] = 4'b0000;
	mem[1528] = 4'b0000;
	mem[1529] = 4'b0000;
	mem[1530] = 4'b0000;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0111;
	mem[1540] = 4'b1100;
	mem[1541] = 4'b1101;
	mem[1542] = 4'b1101;
	mem[1543] = 4'b1101;
	mem[1544] = 4'b1101;
	mem[1545] = 4'b1101;
	mem[1546] = 4'b1101;
	mem[1547] = 4'b1101;
	mem[1548] = 4'b1101;
	mem[1549] = 4'b1101;
	mem[1550] = 4'b1101;
	mem[1551] = 4'b1101;
	mem[1552] = 4'b1101;
	mem[1553] = 4'b1101;
	mem[1554] = 4'b1101;
	mem[1555] = 4'b1101;
	mem[1556] = 4'b1111;
	mem[1557] = 4'b1111;
	mem[1558] = 4'b1111;
	mem[1559] = 4'b1111;
	mem[1560] = 4'b1111;
	mem[1561] = 4'b1111;
	mem[1562] = 4'b1111;
	mem[1563] = 4'b1111;
	mem[1564] = 4'b1111;
	mem[1565] = 4'b1111;
	mem[1566] = 4'b1111;
	mem[1567] = 4'b1111;
	mem[1568] = 4'b1110;
	mem[1569] = 4'b1110;
	mem[1570] = 4'b1111;
	mem[1571] = 4'b1111;
	mem[1572] = 4'b1111;
	mem[1573] = 4'b1111;
	mem[1574] = 4'b1101;
	mem[1575] = 4'b1111;
	mem[1576] = 4'b1111;
	mem[1577] = 4'b1111;
	mem[1578] = 4'b1111;
	mem[1579] = 4'b1111;
	mem[1580] = 4'b1111;
	mem[1581] = 4'b1111;
	mem[1582] = 4'b1111;
	mem[1583] = 4'b1111;
	mem[1584] = 4'b1111;
	mem[1585] = 4'b1111;
	mem[1586] = 4'b1111;
	mem[1587] = 4'b1111;
	mem[1588] = 4'b1111;
	mem[1589] = 4'b1111;
	mem[1590] = 4'b1111;
	mem[1591] = 4'b1111;
	mem[1592] = 4'b1111;
	mem[1593] = 4'b1111;
	mem[1594] = 4'b1111;
	mem[1595] = 4'b1111;
	mem[1596] = 4'b1111;
	mem[1597] = 4'b1111;
	mem[1598] = 4'b1111;
	mem[1599] = 4'b1111;
	mem[1600] = 4'b1111;
	mem[1601] = 4'b1111;
	mem[1602] = 4'b1111;
	mem[1603] = 4'b1111;
	mem[1604] = 4'b1111;
	mem[1605] = 4'b1111;
	mem[1606] = 4'b1111;
	mem[1607] = 4'b1001;
	mem[1608] = 4'b0111;
	mem[1609] = 4'b0111;
	mem[1610] = 4'b0111;
	mem[1611] = 4'b0111;
	mem[1612] = 4'b0110;
	mem[1613] = 4'b0101;
	mem[1614] = 4'b0011;
	mem[1615] = 4'b0001;
	mem[1616] = 4'b0000;
	mem[1617] = 4'b0000;
	mem[1618] = 4'b0000;
	mem[1619] = 4'b0000;
	mem[1620] = 4'b0000;
	mem[1621] = 4'b0000;
	mem[1622] = 4'b0000;
	mem[1623] = 4'b0000;
	mem[1624] = 4'b0001;
	mem[1625] = 4'b0000;
	mem[1626] = 4'b0000;
	mem[1627] = 4'b0000;
	mem[1628] = 4'b0000;
	mem[1629] = 4'b0000;
	mem[1630] = 4'b0001;
	mem[1631] = 4'b0001;
	mem[1632] = 4'b0001;
	mem[1633] = 4'b0000;
	mem[1634] = 4'b0000;
	mem[1635] = 4'b0000;
	mem[1636] = 4'b0000;
	mem[1637] = 4'b0000;
	mem[1638] = 4'b0000;
	mem[1639] = 4'b0000;
	mem[1640] = 4'b0000;
	mem[1641] = 4'b0000;
	mem[1642] = 4'b0000;
	mem[1643] = 4'b0000;
	mem[1644] = 4'b0000;
	mem[1645] = 4'b0000;
	mem[1646] = 4'b0000;
	mem[1647] = 4'b0000;
	mem[1648] = 4'b0000;
	mem[1649] = 4'b0000;
	mem[1650] = 4'b0000;
	mem[1651] = 4'b0000;
	mem[1652] = 4'b0000;
	mem[1653] = 4'b0000;
	mem[1654] = 4'b0000;
	mem[1655] = 4'b0000;
	mem[1656] = 4'b0000;
	mem[1657] = 4'b0000;
	mem[1658] = 4'b0000;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0111;
	mem[1668] = 4'b1100;
	mem[1669] = 4'b1101;
	mem[1670] = 4'b1101;
	mem[1671] = 4'b1101;
	mem[1672] = 4'b1101;
	mem[1673] = 4'b1101;
	mem[1674] = 4'b1101;
	mem[1675] = 4'b1101;
	mem[1676] = 4'b1101;
	mem[1677] = 4'b1101;
	mem[1678] = 4'b1101;
	mem[1679] = 4'b1101;
	mem[1680] = 4'b1101;
	mem[1681] = 4'b1101;
	mem[1682] = 4'b1101;
	mem[1683] = 4'b1101;
	mem[1684] = 4'b1111;
	mem[1685] = 4'b1111;
	mem[1686] = 4'b1111;
	mem[1687] = 4'b1111;
	mem[1688] = 4'b1111;
	mem[1689] = 4'b1111;
	mem[1690] = 4'b1110;
	mem[1691] = 4'b1101;
	mem[1692] = 4'b1101;
	mem[1693] = 4'b1111;
	mem[1694] = 4'b1111;
	mem[1695] = 4'b1111;
	mem[1696] = 4'b1111;
	mem[1697] = 4'b1111;
	mem[1698] = 4'b1111;
	mem[1699] = 4'b1110;
	mem[1700] = 4'b1110;
	mem[1701] = 4'b1101;
	mem[1702] = 4'b1110;
	mem[1703] = 4'b1111;
	mem[1704] = 4'b1111;
	mem[1705] = 4'b1111;
	mem[1706] = 4'b1111;
	mem[1707] = 4'b1111;
	mem[1708] = 4'b1111;
	mem[1709] = 4'b1111;
	mem[1710] = 4'b1111;
	mem[1711] = 4'b1111;
	mem[1712] = 4'b1111;
	mem[1713] = 4'b1111;
	mem[1714] = 4'b1111;
	mem[1715] = 4'b1111;
	mem[1716] = 4'b1111;
	mem[1717] = 4'b1111;
	mem[1718] = 4'b1111;
	mem[1719] = 4'b1111;
	mem[1720] = 4'b1111;
	mem[1721] = 4'b1111;
	mem[1722] = 4'b1111;
	mem[1723] = 4'b1111;
	mem[1724] = 4'b1111;
	mem[1725] = 4'b1111;
	mem[1726] = 4'b1111;
	mem[1727] = 4'b1111;
	mem[1728] = 4'b1111;
	mem[1729] = 4'b1111;
	mem[1730] = 4'b1111;
	mem[1731] = 4'b1111;
	mem[1732] = 4'b1111;
	mem[1733] = 4'b1111;
	mem[1734] = 4'b1111;
	mem[1735] = 4'b1001;
	mem[1736] = 4'b0110;
	mem[1737] = 4'b0101;
	mem[1738] = 4'b0011;
	mem[1739] = 4'b0001;
	mem[1740] = 4'b0000;
	mem[1741] = 4'b0000;
	mem[1742] = 4'b0000;
	mem[1743] = 4'b0000;
	mem[1744] = 4'b0000;
	mem[1745] = 4'b0000;
	mem[1746] = 4'b0000;
	mem[1747] = 4'b0000;
	mem[1748] = 4'b0000;
	mem[1749] = 4'b0000;
	mem[1750] = 4'b0000;
	mem[1751] = 4'b0000;
	mem[1752] = 4'b0001;
	mem[1753] = 4'b0000;
	mem[1754] = 4'b0000;
	mem[1755] = 4'b0000;
	mem[1756] = 4'b0000;
	mem[1757] = 4'b0000;
	mem[1758] = 4'b0001;
	mem[1759] = 4'b0000;
	mem[1760] = 4'b0000;
	mem[1761] = 4'b0000;
	mem[1762] = 4'b0000;
	mem[1763] = 4'b0000;
	mem[1764] = 4'b0000;
	mem[1765] = 4'b0000;
	mem[1766] = 4'b0000;
	mem[1767] = 4'b0000;
	mem[1768] = 4'b0000;
	mem[1769] = 4'b0000;
	mem[1770] = 4'b0000;
	mem[1771] = 4'b0000;
	mem[1772] = 4'b0000;
	mem[1773] = 4'b0000;
	mem[1774] = 4'b0000;
	mem[1775] = 4'b0000;
	mem[1776] = 4'b0000;
	mem[1777] = 4'b0000;
	mem[1778] = 4'b0000;
	mem[1779] = 4'b0000;
	mem[1780] = 4'b0000;
	mem[1781] = 4'b0000;
	mem[1782] = 4'b0000;
	mem[1783] = 4'b0000;
	mem[1784] = 4'b0000;
	mem[1785] = 4'b0000;
	mem[1786] = 4'b0000;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0111;
	mem[1796] = 4'b1100;
	mem[1797] = 4'b1101;
	mem[1798] = 4'b1101;
	mem[1799] = 4'b1101;
	mem[1800] = 4'b1101;
	mem[1801] = 4'b1101;
	mem[1802] = 4'b1101;
	mem[1803] = 4'b1101;
	mem[1804] = 4'b1101;
	mem[1805] = 4'b1101;
	mem[1806] = 4'b1101;
	mem[1807] = 4'b1101;
	mem[1808] = 4'b1101;
	mem[1809] = 4'b1101;
	mem[1810] = 4'b1101;
	mem[1811] = 4'b1101;
	mem[1812] = 4'b1111;
	mem[1813] = 4'b1111;
	mem[1814] = 4'b1111;
	mem[1815] = 4'b1111;
	mem[1816] = 4'b1111;
	mem[1817] = 4'b1110;
	mem[1818] = 4'b1101;
	mem[1819] = 4'b1101;
	mem[1820] = 4'b1101;
	mem[1821] = 4'b1101;
	mem[1822] = 4'b1110;
	mem[1823] = 4'b1111;
	mem[1824] = 4'b1111;
	mem[1825] = 4'b1111;
	mem[1826] = 4'b1101;
	mem[1827] = 4'b1101;
	mem[1828] = 4'b1101;
	mem[1829] = 4'b1110;
	mem[1830] = 4'b1111;
	mem[1831] = 4'b1111;
	mem[1832] = 4'b1111;
	mem[1833] = 4'b1111;
	mem[1834] = 4'b1111;
	mem[1835] = 4'b1111;
	mem[1836] = 4'b1111;
	mem[1837] = 4'b1111;
	mem[1838] = 4'b1111;
	mem[1839] = 4'b1111;
	mem[1840] = 4'b1111;
	mem[1841] = 4'b1111;
	mem[1842] = 4'b1111;
	mem[1843] = 4'b1111;
	mem[1844] = 4'b1111;
	mem[1845] = 4'b1111;
	mem[1846] = 4'b1111;
	mem[1847] = 4'b1111;
	mem[1848] = 4'b1111;
	mem[1849] = 4'b1111;
	mem[1850] = 4'b1111;
	mem[1851] = 4'b1111;
	mem[1852] = 4'b1111;
	mem[1853] = 4'b1111;
	mem[1854] = 4'b1111;
	mem[1855] = 4'b1111;
	mem[1856] = 4'b1111;
	mem[1857] = 4'b1111;
	mem[1858] = 4'b1111;
	mem[1859] = 4'b1111;
	mem[1860] = 4'b1111;
	mem[1861] = 4'b1111;
	mem[1862] = 4'b1111;
	mem[1863] = 4'b0101;
	mem[1864] = 4'b0000;
	mem[1865] = 4'b0000;
	mem[1866] = 4'b0000;
	mem[1867] = 4'b0000;
	mem[1868] = 4'b0000;
	mem[1869] = 4'b0000;
	mem[1870] = 4'b0000;
	mem[1871] = 4'b0000;
	mem[1872] = 4'b0000;
	mem[1873] = 4'b0000;
	mem[1874] = 4'b0000;
	mem[1875] = 4'b0000;
	mem[1876] = 4'b0000;
	mem[1877] = 4'b0000;
	mem[1878] = 4'b0000;
	mem[1879] = 4'b0000;
	mem[1880] = 4'b0000;
	mem[1881] = 4'b0000;
	mem[1882] = 4'b0000;
	mem[1883] = 4'b0000;
	mem[1884] = 4'b0000;
	mem[1885] = 4'b0000;
	mem[1886] = 4'b0001;
	mem[1887] = 4'b0000;
	mem[1888] = 4'b0000;
	mem[1889] = 4'b0000;
	mem[1890] = 4'b0000;
	mem[1891] = 4'b0000;
	mem[1892] = 4'b0000;
	mem[1893] = 4'b0000;
	mem[1894] = 4'b0000;
	mem[1895] = 4'b0000;
	mem[1896] = 4'b0000;
	mem[1897] = 4'b0000;
	mem[1898] = 4'b0000;
	mem[1899] = 4'b0000;
	mem[1900] = 4'b0000;
	mem[1901] = 4'b0000;
	mem[1902] = 4'b0000;
	mem[1903] = 4'b0000;
	mem[1904] = 4'b0000;
	mem[1905] = 4'b0000;
	mem[1906] = 4'b0000;
	mem[1907] = 4'b0000;
	mem[1908] = 4'b0000;
	mem[1909] = 4'b0000;
	mem[1910] = 4'b0000;
	mem[1911] = 4'b0000;
	mem[1912] = 4'b0000;
	mem[1913] = 4'b0000;
	mem[1914] = 4'b0000;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0111;
	mem[1924] = 4'b1100;
	mem[1925] = 4'b1101;
	mem[1926] = 4'b1101;
	mem[1927] = 4'b1101;
	mem[1928] = 4'b1101;
	mem[1929] = 4'b1101;
	mem[1930] = 4'b1101;
	mem[1931] = 4'b1101;
	mem[1932] = 4'b1101;
	mem[1933] = 4'b1101;
	mem[1934] = 4'b1101;
	mem[1935] = 4'b1101;
	mem[1936] = 4'b1101;
	mem[1937] = 4'b1101;
	mem[1938] = 4'b1101;
	mem[1939] = 4'b1110;
	mem[1940] = 4'b1111;
	mem[1941] = 4'b1111;
	mem[1942] = 4'b1111;
	mem[1943] = 4'b1111;
	mem[1944] = 4'b1111;
	mem[1945] = 4'b1101;
	mem[1946] = 4'b1110;
	mem[1947] = 4'b1111;
	mem[1948] = 4'b1110;
	mem[1949] = 4'b1101;
	mem[1950] = 4'b1101;
	mem[1951] = 4'b1110;
	mem[1952] = 4'b1111;
	mem[1953] = 4'b1111;
	mem[1954] = 4'b1111;
	mem[1955] = 4'b1111;
	mem[1956] = 4'b1111;
	mem[1957] = 4'b1111;
	mem[1958] = 4'b1111;
	mem[1959] = 4'b1111;
	mem[1960] = 4'b1111;
	mem[1961] = 4'b1111;
	mem[1962] = 4'b1111;
	mem[1963] = 4'b1111;
	mem[1964] = 4'b1111;
	mem[1965] = 4'b1111;
	mem[1966] = 4'b1111;
	mem[1967] = 4'b1111;
	mem[1968] = 4'b1111;
	mem[1969] = 4'b1111;
	mem[1970] = 4'b1111;
	mem[1971] = 4'b1111;
	mem[1972] = 4'b1111;
	mem[1973] = 4'b1111;
	mem[1974] = 4'b1111;
	mem[1975] = 4'b1111;
	mem[1976] = 4'b1111;
	mem[1977] = 4'b1111;
	mem[1978] = 4'b1111;
	mem[1979] = 4'b1111;
	mem[1980] = 4'b1111;
	mem[1981] = 4'b1111;
	mem[1982] = 4'b1111;
	mem[1983] = 4'b1111;
	mem[1984] = 4'b1110;
	mem[1985] = 4'b1101;
	mem[1986] = 4'b1111;
	mem[1987] = 4'b1111;
	mem[1988] = 4'b1111;
	mem[1989] = 4'b1111;
	mem[1990] = 4'b1111;
	mem[1991] = 4'b0100;
	mem[1992] = 4'b0000;
	mem[1993] = 4'b0000;
	mem[1994] = 4'b0000;
	mem[1995] = 4'b0000;
	mem[1996] = 4'b0000;
	mem[1997] = 4'b0000;
	mem[1998] = 4'b0000;
	mem[1999] = 4'b0000;
	mem[2000] = 4'b0000;
	mem[2001] = 4'b0000;
	mem[2002] = 4'b0000;
	mem[2003] = 4'b0000;
	mem[2004] = 4'b0000;
	mem[2005] = 4'b0000;
	mem[2006] = 4'b0000;
	mem[2007] = 4'b0000;
	mem[2008] = 4'b0000;
	mem[2009] = 4'b0000;
	mem[2010] = 4'b0000;
	mem[2011] = 4'b0000;
	mem[2012] = 4'b0000;
	mem[2013] = 4'b0001;
	mem[2014] = 4'b0000;
	mem[2015] = 4'b0000;
	mem[2016] = 4'b0000;
	mem[2017] = 4'b0000;
	mem[2018] = 4'b0000;
	mem[2019] = 4'b0000;
	mem[2020] = 4'b0000;
	mem[2021] = 4'b0000;
	mem[2022] = 4'b0000;
	mem[2023] = 4'b0000;
	mem[2024] = 4'b0000;
	mem[2025] = 4'b0000;
	mem[2026] = 4'b0000;
	mem[2027] = 4'b0000;
	mem[2028] = 4'b0000;
	mem[2029] = 4'b0000;
	mem[2030] = 4'b0000;
	mem[2031] = 4'b0000;
	mem[2032] = 4'b0000;
	mem[2033] = 4'b0000;
	mem[2034] = 4'b0000;
	mem[2035] = 4'b0000;
	mem[2036] = 4'b0000;
	mem[2037] = 4'b0000;
	mem[2038] = 4'b0000;
	mem[2039] = 4'b0000;
	mem[2040] = 4'b0000;
	mem[2041] = 4'b0000;
	mem[2042] = 4'b0000;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0111;
	mem[2052] = 4'b1100;
	mem[2053] = 4'b1101;
	mem[2054] = 4'b1101;
	mem[2055] = 4'b1101;
	mem[2056] = 4'b1101;
	mem[2057] = 4'b1101;
	mem[2058] = 4'b1101;
	mem[2059] = 4'b1101;
	mem[2060] = 4'b1101;
	mem[2061] = 4'b1101;
	mem[2062] = 4'b1101;
	mem[2063] = 4'b1101;
	mem[2064] = 4'b1101;
	mem[2065] = 4'b1101;
	mem[2066] = 4'b1110;
	mem[2067] = 4'b1110;
	mem[2068] = 4'b1111;
	mem[2069] = 4'b1111;
	mem[2070] = 4'b1111;
	mem[2071] = 4'b1110;
	mem[2072] = 4'b1110;
	mem[2073] = 4'b1110;
	mem[2074] = 4'b1111;
	mem[2075] = 4'b1111;
	mem[2076] = 4'b1111;
	mem[2077] = 4'b1111;
	mem[2078] = 4'b1101;
	mem[2079] = 4'b1101;
	mem[2080] = 4'b1110;
	mem[2081] = 4'b1111;
	mem[2082] = 4'b1111;
	mem[2083] = 4'b1111;
	mem[2084] = 4'b1111;
	mem[2085] = 4'b1111;
	mem[2086] = 4'b1111;
	mem[2087] = 4'b1111;
	mem[2088] = 4'b1111;
	mem[2089] = 4'b1111;
	mem[2090] = 4'b1111;
	mem[2091] = 4'b1111;
	mem[2092] = 4'b1111;
	mem[2093] = 4'b1111;
	mem[2094] = 4'b1111;
	mem[2095] = 4'b1111;
	mem[2096] = 4'b1111;
	mem[2097] = 4'b1111;
	mem[2098] = 4'b1111;
	mem[2099] = 4'b1111;
	mem[2100] = 4'b1111;
	mem[2101] = 4'b1111;
	mem[2102] = 4'b1111;
	mem[2103] = 4'b1111;
	mem[2104] = 4'b1111;
	mem[2105] = 4'b1111;
	mem[2106] = 4'b1111;
	mem[2107] = 4'b1111;
	mem[2108] = 4'b1111;
	mem[2109] = 4'b1111;
	mem[2110] = 4'b1111;
	mem[2111] = 4'b1110;
	mem[2112] = 4'b1101;
	mem[2113] = 4'b1101;
	mem[2114] = 4'b1101;
	mem[2115] = 4'b1111;
	mem[2116] = 4'b1111;
	mem[2117] = 4'b1111;
	mem[2118] = 4'b1111;
	mem[2119] = 4'b0100;
	mem[2120] = 4'b0000;
	mem[2121] = 4'b0000;
	mem[2122] = 4'b0000;
	mem[2123] = 4'b0000;
	mem[2124] = 4'b0000;
	mem[2125] = 4'b0000;
	mem[2126] = 4'b0000;
	mem[2127] = 4'b0000;
	mem[2128] = 4'b0000;
	mem[2129] = 4'b0000;
	mem[2130] = 4'b0000;
	mem[2131] = 4'b0000;
	mem[2132] = 4'b0000;
	mem[2133] = 4'b0000;
	mem[2134] = 4'b0000;
	mem[2135] = 4'b0000;
	mem[2136] = 4'b0000;
	mem[2137] = 4'b0000;
	mem[2138] = 4'b0000;
	mem[2139] = 4'b0000;
	mem[2140] = 4'b0001;
	mem[2141] = 4'b0001;
	mem[2142] = 4'b0000;
	mem[2143] = 4'b0000;
	mem[2144] = 4'b0000;
	mem[2145] = 4'b0000;
	mem[2146] = 4'b0000;
	mem[2147] = 4'b0000;
	mem[2148] = 4'b0000;
	mem[2149] = 4'b0000;
	mem[2150] = 4'b0000;
	mem[2151] = 4'b0000;
	mem[2152] = 4'b0000;
	mem[2153] = 4'b0000;
	mem[2154] = 4'b0000;
	mem[2155] = 4'b0000;
	mem[2156] = 4'b0000;
	mem[2157] = 4'b0000;
	mem[2158] = 4'b0000;
	mem[2159] = 4'b0000;
	mem[2160] = 4'b0000;
	mem[2161] = 4'b0000;
	mem[2162] = 4'b0000;
	mem[2163] = 4'b0000;
	mem[2164] = 4'b0000;
	mem[2165] = 4'b0000;
	mem[2166] = 4'b0000;
	mem[2167] = 4'b0000;
	mem[2168] = 4'b0000;
	mem[2169] = 4'b0000;
	mem[2170] = 4'b0000;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0111;
	mem[2180] = 4'b1100;
	mem[2181] = 4'b1101;
	mem[2182] = 4'b1101;
	mem[2183] = 4'b1101;
	mem[2184] = 4'b1101;
	mem[2185] = 4'b1101;
	mem[2186] = 4'b1101;
	mem[2187] = 4'b1101;
	mem[2188] = 4'b1101;
	mem[2189] = 4'b1101;
	mem[2190] = 4'b1101;
	mem[2191] = 4'b1101;
	mem[2192] = 4'b1110;
	mem[2193] = 4'b1110;
	mem[2194] = 4'b1110;
	mem[2195] = 4'b1110;
	mem[2196] = 4'b1111;
	mem[2197] = 4'b1111;
	mem[2198] = 4'b1111;
	mem[2199] = 4'b1101;
	mem[2200] = 4'b1101;
	mem[2201] = 4'b1101;
	mem[2202] = 4'b1111;
	mem[2203] = 4'b1111;
	mem[2204] = 4'b1111;
	mem[2205] = 4'b1111;
	mem[2206] = 4'b1111;
	mem[2207] = 4'b1101;
	mem[2208] = 4'b1101;
	mem[2209] = 4'b1110;
	mem[2210] = 4'b1111;
	mem[2211] = 4'b1111;
	mem[2212] = 4'b1111;
	mem[2213] = 4'b1111;
	mem[2214] = 4'b1111;
	mem[2215] = 4'b1111;
	mem[2216] = 4'b1111;
	mem[2217] = 4'b1111;
	mem[2218] = 4'b1111;
	mem[2219] = 4'b1111;
	mem[2220] = 4'b1111;
	mem[2221] = 4'b1111;
	mem[2222] = 4'b1111;
	mem[2223] = 4'b1111;
	mem[2224] = 4'b1111;
	mem[2225] = 4'b1111;
	mem[2226] = 4'b1111;
	mem[2227] = 4'b1111;
	mem[2228] = 4'b1111;
	mem[2229] = 4'b1111;
	mem[2230] = 4'b1111;
	mem[2231] = 4'b1111;
	mem[2232] = 4'b1111;
	mem[2233] = 4'b1111;
	mem[2234] = 4'b1111;
	mem[2235] = 4'b1111;
	mem[2236] = 4'b1111;
	mem[2237] = 4'b1111;
	mem[2238] = 4'b1111;
	mem[2239] = 4'b1101;
	mem[2240] = 4'b1101;
	mem[2241] = 4'b1101;
	mem[2242] = 4'b1101;
	mem[2243] = 4'b1101;
	mem[2244] = 4'b1111;
	mem[2245] = 4'b1111;
	mem[2246] = 4'b1111;
	mem[2247] = 4'b0100;
	mem[2248] = 4'b0000;
	mem[2249] = 4'b0000;
	mem[2250] = 4'b0000;
	mem[2251] = 4'b0000;
	mem[2252] = 4'b0000;
	mem[2253] = 4'b0000;
	mem[2254] = 4'b0000;
	mem[2255] = 4'b0000;
	mem[2256] = 4'b0000;
	mem[2257] = 4'b0000;
	mem[2258] = 4'b0000;
	mem[2259] = 4'b0000;
	mem[2260] = 4'b0000;
	mem[2261] = 4'b0000;
	mem[2262] = 4'b0000;
	mem[2263] = 4'b0000;
	mem[2264] = 4'b0000;
	mem[2265] = 4'b0000;
	mem[2266] = 4'b0000;
	mem[2267] = 4'b0001;
	mem[2268] = 4'b0001;
	mem[2269] = 4'b0000;
	mem[2270] = 4'b0000;
	mem[2271] = 4'b0000;
	mem[2272] = 4'b0000;
	mem[2273] = 4'b0000;
	mem[2274] = 4'b0000;
	mem[2275] = 4'b0000;
	mem[2276] = 4'b0000;
	mem[2277] = 4'b0000;
	mem[2278] = 4'b0000;
	mem[2279] = 4'b0000;
	mem[2280] = 4'b0000;
	mem[2281] = 4'b0000;
	mem[2282] = 4'b0000;
	mem[2283] = 4'b0000;
	mem[2284] = 4'b0000;
	mem[2285] = 4'b0000;
	mem[2286] = 4'b0000;
	mem[2287] = 4'b0000;
	mem[2288] = 4'b0000;
	mem[2289] = 4'b0000;
	mem[2290] = 4'b0000;
	mem[2291] = 4'b0000;
	mem[2292] = 4'b0000;
	mem[2293] = 4'b0000;
	mem[2294] = 4'b0000;
	mem[2295] = 4'b0000;
	mem[2296] = 4'b0000;
	mem[2297] = 4'b0000;
	mem[2298] = 4'b0000;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0111;
	mem[2308] = 4'b1100;
	mem[2309] = 4'b1101;
	mem[2310] = 4'b1101;
	mem[2311] = 4'b1101;
	mem[2312] = 4'b1101;
	mem[2313] = 4'b1101;
	mem[2314] = 4'b1101;
	mem[2315] = 4'b1101;
	mem[2316] = 4'b1101;
	mem[2317] = 4'b1101;
	mem[2318] = 4'b1110;
	mem[2319] = 4'b1110;
	mem[2320] = 4'b1110;
	mem[2321] = 4'b1110;
	mem[2322] = 4'b1110;
	mem[2323] = 4'b1110;
	mem[2324] = 4'b1111;
	mem[2325] = 4'b1111;
	mem[2326] = 4'b1111;
	mem[2327] = 4'b1111;
	mem[2328] = 4'b1101;
	mem[2329] = 4'b1101;
	mem[2330] = 4'b1110;
	mem[2331] = 4'b1111;
	mem[2332] = 4'b1111;
	mem[2333] = 4'b1111;
	mem[2334] = 4'b1111;
	mem[2335] = 4'b1111;
	mem[2336] = 4'b1101;
	mem[2337] = 4'b1110;
	mem[2338] = 4'b1111;
	mem[2339] = 4'b1111;
	mem[2340] = 4'b1111;
	mem[2341] = 4'b1111;
	mem[2342] = 4'b1111;
	mem[2343] = 4'b1111;
	mem[2344] = 4'b1111;
	mem[2345] = 4'b1111;
	mem[2346] = 4'b1111;
	mem[2347] = 4'b1111;
	mem[2348] = 4'b1111;
	mem[2349] = 4'b1111;
	mem[2350] = 4'b1111;
	mem[2351] = 4'b1111;
	mem[2352] = 4'b1111;
	mem[2353] = 4'b1111;
	mem[2354] = 4'b1111;
	mem[2355] = 4'b1111;
	mem[2356] = 4'b1111;
	mem[2357] = 4'b1111;
	mem[2358] = 4'b1111;
	mem[2359] = 4'b1111;
	mem[2360] = 4'b1111;
	mem[2361] = 4'b1111;
	mem[2362] = 4'b1111;
	mem[2363] = 4'b1111;
	mem[2364] = 4'b1111;
	mem[2365] = 4'b1111;
	mem[2366] = 4'b1111;
	mem[2367] = 4'b1111;
	mem[2368] = 4'b1101;
	mem[2369] = 4'b1101;
	mem[2370] = 4'b1101;
	mem[2371] = 4'b1101;
	mem[2372] = 4'b1101;
	mem[2373] = 4'b1111;
	mem[2374] = 4'b1111;
	mem[2375] = 4'b0100;
	mem[2376] = 4'b0000;
	mem[2377] = 4'b0000;
	mem[2378] = 4'b0000;
	mem[2379] = 4'b0000;
	mem[2380] = 4'b0000;
	mem[2381] = 4'b0000;
	mem[2382] = 4'b0000;
	mem[2383] = 4'b0000;
	mem[2384] = 4'b0000;
	mem[2385] = 4'b0000;
	mem[2386] = 4'b0000;
	mem[2387] = 4'b0000;
	mem[2388] = 4'b0000;
	mem[2389] = 4'b0000;
	mem[2390] = 4'b0000;
	mem[2391] = 4'b0000;
	mem[2392] = 4'b0001;
	mem[2393] = 4'b0001;
	mem[2394] = 4'b0001;
	mem[2395] = 4'b0000;
	mem[2396] = 4'b0000;
	mem[2397] = 4'b0000;
	mem[2398] = 4'b0000;
	mem[2399] = 4'b0000;
	mem[2400] = 4'b0000;
	mem[2401] = 4'b0000;
	mem[2402] = 4'b0000;
	mem[2403] = 4'b0000;
	mem[2404] = 4'b0000;
	mem[2405] = 4'b0000;
	mem[2406] = 4'b0000;
	mem[2407] = 4'b0000;
	mem[2408] = 4'b0000;
	mem[2409] = 4'b0000;
	mem[2410] = 4'b0000;
	mem[2411] = 4'b0000;
	mem[2412] = 4'b0000;
	mem[2413] = 4'b0000;
	mem[2414] = 4'b0000;
	mem[2415] = 4'b0000;
	mem[2416] = 4'b0000;
	mem[2417] = 4'b0000;
	mem[2418] = 4'b0000;
	mem[2419] = 4'b0000;
	mem[2420] = 4'b0000;
	mem[2421] = 4'b0000;
	mem[2422] = 4'b0000;
	mem[2423] = 4'b0000;
	mem[2424] = 4'b0000;
	mem[2425] = 4'b0000;
	mem[2426] = 4'b0000;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0111;
	mem[2436] = 4'b1100;
	mem[2437] = 4'b1101;
	mem[2438] = 4'b1101;
	mem[2439] = 4'b1101;
	mem[2440] = 4'b1101;
	mem[2441] = 4'b1101;
	mem[2442] = 4'b1101;
	mem[2443] = 4'b1101;
	mem[2444] = 4'b1110;
	mem[2445] = 4'b1110;
	mem[2446] = 4'b1110;
	mem[2447] = 4'b1110;
	mem[2448] = 4'b1110;
	mem[2449] = 4'b1110;
	mem[2450] = 4'b1110;
	mem[2451] = 4'b1110;
	mem[2452] = 4'b1111;
	mem[2453] = 4'b1111;
	mem[2454] = 4'b1111;
	mem[2455] = 4'b1111;
	mem[2456] = 4'b1111;
	mem[2457] = 4'b1101;
	mem[2458] = 4'b1101;
	mem[2459] = 4'b1110;
	mem[2460] = 4'b1111;
	mem[2461] = 4'b1111;
	mem[2462] = 4'b1111;
	mem[2463] = 4'b1111;
	mem[2464] = 4'b1111;
	mem[2465] = 4'b1111;
	mem[2466] = 4'b1111;
	mem[2467] = 4'b1111;
	mem[2468] = 4'b1111;
	mem[2469] = 4'b1111;
	mem[2470] = 4'b1111;
	mem[2471] = 4'b1111;
	mem[2472] = 4'b1111;
	mem[2473] = 4'b1111;
	mem[2474] = 4'b1111;
	mem[2475] = 4'b1111;
	mem[2476] = 4'b1111;
	mem[2477] = 4'b1111;
	mem[2478] = 4'b1111;
	mem[2479] = 4'b1111;
	mem[2480] = 4'b1111;
	mem[2481] = 4'b1111;
	mem[2482] = 4'b1111;
	mem[2483] = 4'b1111;
	mem[2484] = 4'b1111;
	mem[2485] = 4'b1111;
	mem[2486] = 4'b1111;
	mem[2487] = 4'b1111;
	mem[2488] = 4'b1111;
	mem[2489] = 4'b1111;
	mem[2490] = 4'b1111;
	mem[2491] = 4'b1111;
	mem[2492] = 4'b1111;
	mem[2493] = 4'b1111;
	mem[2494] = 4'b1111;
	mem[2495] = 4'b1111;
	mem[2496] = 4'b1111;
	mem[2497] = 4'b1101;
	mem[2498] = 4'b1101;
	mem[2499] = 4'b1101;
	mem[2500] = 4'b1101;
	mem[2501] = 4'b1101;
	mem[2502] = 4'b1111;
	mem[2503] = 4'b0100;
	mem[2504] = 4'b0000;
	mem[2505] = 4'b0000;
	mem[2506] = 4'b0000;
	mem[2507] = 4'b0000;
	mem[2508] = 4'b0000;
	mem[2509] = 4'b0000;
	mem[2510] = 4'b0000;
	mem[2511] = 4'b0000;
	mem[2512] = 4'b0000;
	mem[2513] = 4'b0000;
	mem[2514] = 4'b0000;
	mem[2515] = 4'b0000;
	mem[2516] = 4'b0000;
	mem[2517] = 4'b0000;
	mem[2518] = 4'b0000;
	mem[2519] = 4'b0000;
	mem[2520] = 4'b0000;
	mem[2521] = 4'b0000;
	mem[2522] = 4'b0000;
	mem[2523] = 4'b0000;
	mem[2524] = 4'b0000;
	mem[2525] = 4'b0000;
	mem[2526] = 4'b0000;
	mem[2527] = 4'b0000;
	mem[2528] = 4'b0000;
	mem[2529] = 4'b0000;
	mem[2530] = 4'b0000;
	mem[2531] = 4'b0000;
	mem[2532] = 4'b0000;
	mem[2533] = 4'b0000;
	mem[2534] = 4'b0000;
	mem[2535] = 4'b0000;
	mem[2536] = 4'b0000;
	mem[2537] = 4'b0000;
	mem[2538] = 4'b0000;
	mem[2539] = 4'b0000;
	mem[2540] = 4'b0000;
	mem[2541] = 4'b0000;
	mem[2542] = 4'b0000;
	mem[2543] = 4'b0000;
	mem[2544] = 4'b0000;
	mem[2545] = 4'b0000;
	mem[2546] = 4'b0000;
	mem[2547] = 4'b0000;
	mem[2548] = 4'b0000;
	mem[2549] = 4'b0000;
	mem[2550] = 4'b0000;
	mem[2551] = 4'b0000;
	mem[2552] = 4'b0000;
	mem[2553] = 4'b0000;
	mem[2554] = 4'b0000;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b0111;
	mem[2564] = 4'b1100;
	mem[2565] = 4'b1101;
	mem[2566] = 4'b1101;
	mem[2567] = 4'b1101;
	mem[2568] = 4'b1101;
	mem[2569] = 4'b1101;
	mem[2570] = 4'b1110;
	mem[2571] = 4'b1110;
	mem[2572] = 4'b1110;
	mem[2573] = 4'b1110;
	mem[2574] = 4'b1110;
	mem[2575] = 4'b1110;
	mem[2576] = 4'b1110;
	mem[2577] = 4'b1110;
	mem[2578] = 4'b1101;
	mem[2579] = 4'b1101;
	mem[2580] = 4'b1110;
	mem[2581] = 4'b1110;
	mem[2582] = 4'b1111;
	mem[2583] = 4'b1111;
	mem[2584] = 4'b1111;
	mem[2585] = 4'b1111;
	mem[2586] = 4'b1101;
	mem[2587] = 4'b1101;
	mem[2588] = 4'b1110;
	mem[2589] = 4'b1111;
	mem[2590] = 4'b1111;
	mem[2591] = 4'b1111;
	mem[2592] = 4'b1111;
	mem[2593] = 4'b1111;
	mem[2594] = 4'b1111;
	mem[2595] = 4'b1111;
	mem[2596] = 4'b1111;
	mem[2597] = 4'b1111;
	mem[2598] = 4'b1111;
	mem[2599] = 4'b1111;
	mem[2600] = 4'b1111;
	mem[2601] = 4'b1111;
	mem[2602] = 4'b1111;
	mem[2603] = 4'b1111;
	mem[2604] = 4'b1111;
	mem[2605] = 4'b1111;
	mem[2606] = 4'b1111;
	mem[2607] = 4'b1111;
	mem[2608] = 4'b1111;
	mem[2609] = 4'b1111;
	mem[2610] = 4'b1111;
	mem[2611] = 4'b1111;
	mem[2612] = 4'b1111;
	mem[2613] = 4'b1111;
	mem[2614] = 4'b1111;
	mem[2615] = 4'b1111;
	mem[2616] = 4'b1111;
	mem[2617] = 4'b1111;
	mem[2618] = 4'b1111;
	mem[2619] = 4'b1111;
	mem[2620] = 4'b1111;
	mem[2621] = 4'b1111;
	mem[2622] = 4'b1111;
	mem[2623] = 4'b1111;
	mem[2624] = 4'b1111;
	mem[2625] = 4'b1111;
	mem[2626] = 4'b1101;
	mem[2627] = 4'b1101;
	mem[2628] = 4'b1101;
	mem[2629] = 4'b1101;
	mem[2630] = 4'b1101;
	mem[2631] = 4'b0100;
	mem[2632] = 4'b0000;
	mem[2633] = 4'b0000;
	mem[2634] = 4'b0000;
	mem[2635] = 4'b0000;
	mem[2636] = 4'b0000;
	mem[2637] = 4'b0000;
	mem[2638] = 4'b0000;
	mem[2639] = 4'b0000;
	mem[2640] = 4'b0000;
	mem[2641] = 4'b0000;
	mem[2642] = 4'b0000;
	mem[2643] = 4'b0000;
	mem[2644] = 4'b0000;
	mem[2645] = 4'b0000;
	mem[2646] = 4'b0000;
	mem[2647] = 4'b0000;
	mem[2648] = 4'b0000;
	mem[2649] = 4'b0000;
	mem[2650] = 4'b0000;
	mem[2651] = 4'b0000;
	mem[2652] = 4'b0000;
	mem[2653] = 4'b0000;
	mem[2654] = 4'b0000;
	mem[2655] = 4'b0000;
	mem[2656] = 4'b0000;
	mem[2657] = 4'b0000;
	mem[2658] = 4'b0000;
	mem[2659] = 4'b0000;
	mem[2660] = 4'b0000;
	mem[2661] = 4'b0000;
	mem[2662] = 4'b0000;
	mem[2663] = 4'b0000;
	mem[2664] = 4'b0000;
	mem[2665] = 4'b0000;
	mem[2666] = 4'b0000;
	mem[2667] = 4'b0000;
	mem[2668] = 4'b0000;
	mem[2669] = 4'b0000;
	mem[2670] = 4'b0000;
	mem[2671] = 4'b0000;
	mem[2672] = 4'b0000;
	mem[2673] = 4'b0000;
	mem[2674] = 4'b0000;
	mem[2675] = 4'b0000;
	mem[2676] = 4'b0000;
	mem[2677] = 4'b0000;
	mem[2678] = 4'b0000;
	mem[2679] = 4'b0000;
	mem[2680] = 4'b0000;
	mem[2681] = 4'b0000;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b0111;
	mem[2692] = 4'b1100;
	mem[2693] = 4'b1101;
	mem[2694] = 4'b1101;
	mem[2695] = 4'b1101;
	mem[2696] = 4'b1110;
	mem[2697] = 4'b1110;
	mem[2698] = 4'b1110;
	mem[2699] = 4'b1110;
	mem[2700] = 4'b1110;
	mem[2701] = 4'b1110;
	mem[2702] = 4'b1110;
	mem[2703] = 4'b1110;
	mem[2704] = 4'b1110;
	mem[2705] = 4'b1101;
	mem[2706] = 4'b1100;
	mem[2707] = 4'b1100;
	mem[2708] = 4'b1101;
	mem[2709] = 4'b1101;
	mem[2710] = 4'b1101;
	mem[2711] = 4'b1110;
	mem[2712] = 4'b1111;
	mem[2713] = 4'b1111;
	mem[2714] = 4'b1111;
	mem[2715] = 4'b1101;
	mem[2716] = 4'b1101;
	mem[2717] = 4'b1110;
	mem[2718] = 4'b1111;
	mem[2719] = 4'b1111;
	mem[2720] = 4'b1111;
	mem[2721] = 4'b1111;
	mem[2722] = 4'b1111;
	mem[2723] = 4'b1111;
	mem[2724] = 4'b1111;
	mem[2725] = 4'b1111;
	mem[2726] = 4'b1111;
	mem[2727] = 4'b1111;
	mem[2728] = 4'b1111;
	mem[2729] = 4'b1111;
	mem[2730] = 4'b1111;
	mem[2731] = 4'b1111;
	mem[2732] = 4'b1111;
	mem[2733] = 4'b1111;
	mem[2734] = 4'b1111;
	mem[2735] = 4'b1111;
	mem[2736] = 4'b1111;
	mem[2737] = 4'b1111;
	mem[2738] = 4'b1111;
	mem[2739] = 4'b1111;
	mem[2740] = 4'b1111;
	mem[2741] = 4'b1111;
	mem[2742] = 4'b1111;
	mem[2743] = 4'b1111;
	mem[2744] = 4'b1111;
	mem[2745] = 4'b1111;
	mem[2746] = 4'b1111;
	mem[2747] = 4'b1111;
	mem[2748] = 4'b1111;
	mem[2749] = 4'b1111;
	mem[2750] = 4'b1111;
	mem[2751] = 4'b1111;
	mem[2752] = 4'b1111;
	mem[2753] = 4'b1111;
	mem[2754] = 4'b1111;
	mem[2755] = 4'b1101;
	mem[2756] = 4'b1101;
	mem[2757] = 4'b1101;
	mem[2758] = 4'b1101;
	mem[2759] = 4'b0011;
	mem[2760] = 4'b0000;
	mem[2761] = 4'b0000;
	mem[2762] = 4'b0000;
	mem[2763] = 4'b0000;
	mem[2764] = 4'b0000;
	mem[2765] = 4'b0000;
	mem[2766] = 4'b0000;
	mem[2767] = 4'b0000;
	mem[2768] = 4'b0000;
	mem[2769] = 4'b0000;
	mem[2770] = 4'b0000;
	mem[2771] = 4'b0000;
	mem[2772] = 4'b0000;
	mem[2773] = 4'b0000;
	mem[2774] = 4'b0000;
	mem[2775] = 4'b0000;
	mem[2776] = 4'b0000;
	mem[2777] = 4'b0000;
	mem[2778] = 4'b0000;
	mem[2779] = 4'b0000;
	mem[2780] = 4'b0000;
	mem[2781] = 4'b0000;
	mem[2782] = 4'b0000;
	mem[2783] = 4'b0000;
	mem[2784] = 4'b0000;
	mem[2785] = 4'b0000;
	mem[2786] = 4'b0000;
	mem[2787] = 4'b0000;
	mem[2788] = 4'b0000;
	mem[2789] = 4'b0000;
	mem[2790] = 4'b0000;
	mem[2791] = 4'b0000;
	mem[2792] = 4'b0000;
	mem[2793] = 4'b0000;
	mem[2794] = 4'b0000;
	mem[2795] = 4'b0000;
	mem[2796] = 4'b0000;
	mem[2797] = 4'b0000;
	mem[2798] = 4'b0000;
	mem[2799] = 4'b0000;
	mem[2800] = 4'b0000;
	mem[2801] = 4'b0000;
	mem[2802] = 4'b0000;
	mem[2803] = 4'b0000;
	mem[2804] = 4'b0000;
	mem[2805] = 4'b0000;
	mem[2806] = 4'b0000;
	mem[2807] = 4'b0000;
	mem[2808] = 4'b0000;
	mem[2809] = 4'b0000;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b0111;
	mem[2820] = 4'b1100;
	mem[2821] = 4'b1101;
	mem[2822] = 4'b1101;
	mem[2823] = 4'b1110;
	mem[2824] = 4'b1110;
	mem[2825] = 4'b1110;
	mem[2826] = 4'b1110;
	mem[2827] = 4'b1110;
	mem[2828] = 4'b1110;
	mem[2829] = 4'b1110;
	mem[2830] = 4'b1110;
	mem[2831] = 4'b1110;
	mem[2832] = 4'b1101;
	mem[2833] = 4'b1100;
	mem[2834] = 4'b1100;
	mem[2835] = 4'b1101;
	mem[2836] = 4'b1111;
	mem[2837] = 4'b1111;
	mem[2838] = 4'b1101;
	mem[2839] = 4'b1101;
	mem[2840] = 4'b1110;
	mem[2841] = 4'b1111;
	mem[2842] = 4'b1111;
	mem[2843] = 4'b1111;
	mem[2844] = 4'b1101;
	mem[2845] = 4'b1110;
	mem[2846] = 4'b1111;
	mem[2847] = 4'b1111;
	mem[2848] = 4'b1111;
	mem[2849] = 4'b1111;
	mem[2850] = 4'b1111;
	mem[2851] = 4'b1111;
	mem[2852] = 4'b1111;
	mem[2853] = 4'b1111;
	mem[2854] = 4'b1111;
	mem[2855] = 4'b1111;
	mem[2856] = 4'b1111;
	mem[2857] = 4'b1111;
	mem[2858] = 4'b1111;
	mem[2859] = 4'b1111;
	mem[2860] = 4'b1111;
	mem[2861] = 4'b1111;
	mem[2862] = 4'b1111;
	mem[2863] = 4'b1111;
	mem[2864] = 4'b1111;
	mem[2865] = 4'b1111;
	mem[2866] = 4'b1111;
	mem[2867] = 4'b1111;
	mem[2868] = 4'b1111;
	mem[2869] = 4'b1111;
	mem[2870] = 4'b1111;
	mem[2871] = 4'b1111;
	mem[2872] = 4'b1111;
	mem[2873] = 4'b1111;
	mem[2874] = 4'b1111;
	mem[2875] = 4'b1111;
	mem[2876] = 4'b1111;
	mem[2877] = 4'b1111;
	mem[2878] = 4'b1111;
	mem[2879] = 4'b1111;
	mem[2880] = 4'b1111;
	mem[2881] = 4'b1111;
	mem[2882] = 4'b1111;
	mem[2883] = 4'b1111;
	mem[2884] = 4'b1101;
	mem[2885] = 4'b1101;
	mem[2886] = 4'b1101;
	mem[2887] = 4'b0011;
	mem[2888] = 4'b0000;
	mem[2889] = 4'b0000;
	mem[2890] = 4'b0000;
	mem[2891] = 4'b0000;
	mem[2892] = 4'b0000;
	mem[2893] = 4'b0000;
	mem[2894] = 4'b0000;
	mem[2895] = 4'b0000;
	mem[2896] = 4'b0000;
	mem[2897] = 4'b0000;
	mem[2898] = 4'b0000;
	mem[2899] = 4'b0000;
	mem[2900] = 4'b0000;
	mem[2901] = 4'b0000;
	mem[2902] = 4'b0001;
	mem[2903] = 4'b0001;
	mem[2904] = 4'b0000;
	mem[2905] = 4'b0000;
	mem[2906] = 4'b0000;
	mem[2907] = 4'b0000;
	mem[2908] = 4'b0000;
	mem[2909] = 4'b0000;
	mem[2910] = 4'b0000;
	mem[2911] = 4'b0000;
	mem[2912] = 4'b0000;
	mem[2913] = 4'b0000;
	mem[2914] = 4'b0000;
	mem[2915] = 4'b0000;
	mem[2916] = 4'b0000;
	mem[2917] = 4'b0000;
	mem[2918] = 4'b0000;
	mem[2919] = 4'b0000;
	mem[2920] = 4'b0000;
	mem[2921] = 4'b0000;
	mem[2922] = 4'b0000;
	mem[2923] = 4'b0000;
	mem[2924] = 4'b0000;
	mem[2925] = 4'b0000;
	mem[2926] = 4'b0000;
	mem[2927] = 4'b0000;
	mem[2928] = 4'b0000;
	mem[2929] = 4'b0000;
	mem[2930] = 4'b0000;
	mem[2931] = 4'b0000;
	mem[2932] = 4'b0000;
	mem[2933] = 4'b0000;
	mem[2934] = 4'b0000;
	mem[2935] = 4'b0000;
	mem[2936] = 4'b0000;
	mem[2937] = 4'b0000;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b0111;
	mem[2948] = 4'b1100;
	mem[2949] = 4'b1101;
	mem[2950] = 4'b1110;
	mem[2951] = 4'b1110;
	mem[2952] = 4'b1110;
	mem[2953] = 4'b1110;
	mem[2954] = 4'b1110;
	mem[2955] = 4'b1110;
	mem[2956] = 4'b1110;
	mem[2957] = 4'b1110;
	mem[2958] = 4'b1110;
	mem[2959] = 4'b1110;
	mem[2960] = 4'b1101;
	mem[2961] = 4'b1100;
	mem[2962] = 4'b1100;
	mem[2963] = 4'b1110;
	mem[2964] = 4'b1111;
	mem[2965] = 4'b1111;
	mem[2966] = 4'b1111;
	mem[2967] = 4'b1101;
	mem[2968] = 4'b1101;
	mem[2969] = 4'b1111;
	mem[2970] = 4'b1111;
	mem[2971] = 4'b1111;
	mem[2972] = 4'b1111;
	mem[2973] = 4'b1111;
	mem[2974] = 4'b1111;
	mem[2975] = 4'b1111;
	mem[2976] = 4'b1111;
	mem[2977] = 4'b1111;
	mem[2978] = 4'b1111;
	mem[2979] = 4'b1111;
	mem[2980] = 4'b1111;
	mem[2981] = 4'b1111;
	mem[2982] = 4'b1111;
	mem[2983] = 4'b1111;
	mem[2984] = 4'b1111;
	mem[2985] = 4'b1111;
	mem[2986] = 4'b1111;
	mem[2987] = 4'b1111;
	mem[2988] = 4'b1111;
	mem[2989] = 4'b1111;
	mem[2990] = 4'b1111;
	mem[2991] = 4'b1111;
	mem[2992] = 4'b1111;
	mem[2993] = 4'b1111;
	mem[2994] = 4'b1111;
	mem[2995] = 4'b1111;
	mem[2996] = 4'b1111;
	mem[2997] = 4'b1111;
	mem[2998] = 4'b1111;
	mem[2999] = 4'b1111;
	mem[3000] = 4'b1111;
	mem[3001] = 4'b1111;
	mem[3002] = 4'b1111;
	mem[3003] = 4'b1111;
	mem[3004] = 4'b1111;
	mem[3005] = 4'b1111;
	mem[3006] = 4'b1111;
	mem[3007] = 4'b1111;
	mem[3008] = 4'b1111;
	mem[3009] = 4'b1111;
	mem[3010] = 4'b1111;
	mem[3011] = 4'b1111;
	mem[3012] = 4'b1111;
	mem[3013] = 4'b1101;
	mem[3014] = 4'b1101;
	mem[3015] = 4'b0011;
	mem[3016] = 4'b0000;
	mem[3017] = 4'b0000;
	mem[3018] = 4'b0000;
	mem[3019] = 4'b0000;
	mem[3020] = 4'b0000;
	mem[3021] = 4'b0000;
	mem[3022] = 4'b0000;
	mem[3023] = 4'b0000;
	mem[3024] = 4'b0000;
	mem[3025] = 4'b0000;
	mem[3026] = 4'b0000;
	mem[3027] = 4'b0000;
	mem[3028] = 4'b0000;
	mem[3029] = 4'b0001;
	mem[3030] = 4'b0001;
	mem[3031] = 4'b0000;
	mem[3032] = 4'b0000;
	mem[3033] = 4'b0000;
	mem[3034] = 4'b0000;
	mem[3035] = 4'b0000;
	mem[3036] = 4'b0000;
	mem[3037] = 4'b0000;
	mem[3038] = 4'b0000;
	mem[3039] = 4'b0000;
	mem[3040] = 4'b0000;
	mem[3041] = 4'b0000;
	mem[3042] = 4'b0000;
	mem[3043] = 4'b0000;
	mem[3044] = 4'b0000;
	mem[3045] = 4'b0000;
	mem[3046] = 4'b0000;
	mem[3047] = 4'b0000;
	mem[3048] = 4'b0000;
	mem[3049] = 4'b0000;
	mem[3050] = 4'b0000;
	mem[3051] = 4'b0000;
	mem[3052] = 4'b0000;
	mem[3053] = 4'b0000;
	mem[3054] = 4'b0000;
	mem[3055] = 4'b0000;
	mem[3056] = 4'b0000;
	mem[3057] = 4'b0000;
	mem[3058] = 4'b0000;
	mem[3059] = 4'b0000;
	mem[3060] = 4'b0000;
	mem[3061] = 4'b0000;
	mem[3062] = 4'b0000;
	mem[3063] = 4'b0000;
	mem[3064] = 4'b0000;
	mem[3065] = 4'b0000;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b0111;
	mem[3076] = 4'b1100;
	mem[3077] = 4'b1101;
	mem[3078] = 4'b1110;
	mem[3079] = 4'b1110;
	mem[3080] = 4'b1110;
	mem[3081] = 4'b1110;
	mem[3082] = 4'b1110;
	mem[3083] = 4'b1110;
	mem[3084] = 4'b1110;
	mem[3085] = 4'b1110;
	mem[3086] = 4'b1110;
	mem[3087] = 4'b1110;
	mem[3088] = 4'b1101;
	mem[3089] = 4'b1100;
	mem[3090] = 4'b1101;
	mem[3091] = 4'b1110;
	mem[3092] = 4'b1111;
	mem[3093] = 4'b1111;
	mem[3094] = 4'b1111;
	mem[3095] = 4'b1111;
	mem[3096] = 4'b1101;
	mem[3097] = 4'b1110;
	mem[3098] = 4'b1111;
	mem[3099] = 4'b1111;
	mem[3100] = 4'b1111;
	mem[3101] = 4'b1111;
	mem[3102] = 4'b1111;
	mem[3103] = 4'b1111;
	mem[3104] = 4'b1111;
	mem[3105] = 4'b1111;
	mem[3106] = 4'b1111;
	mem[3107] = 4'b1111;
	mem[3108] = 4'b1111;
	mem[3109] = 4'b1111;
	mem[3110] = 4'b1111;
	mem[3111] = 4'b1111;
	mem[3112] = 4'b1111;
	mem[3113] = 4'b1111;
	mem[3114] = 4'b1111;
	mem[3115] = 4'b1111;
	mem[3116] = 4'b1111;
	mem[3117] = 4'b1111;
	mem[3118] = 4'b1111;
	mem[3119] = 4'b1111;
	mem[3120] = 4'b1111;
	mem[3121] = 4'b1111;
	mem[3122] = 4'b1111;
	mem[3123] = 4'b1111;
	mem[3124] = 4'b1111;
	mem[3125] = 4'b1111;
	mem[3126] = 4'b1111;
	mem[3127] = 4'b1111;
	mem[3128] = 4'b1111;
	mem[3129] = 4'b1111;
	mem[3130] = 4'b1111;
	mem[3131] = 4'b1111;
	mem[3132] = 4'b1111;
	mem[3133] = 4'b1111;
	mem[3134] = 4'b1111;
	mem[3135] = 4'b1111;
	mem[3136] = 4'b1111;
	mem[3137] = 4'b1111;
	mem[3138] = 4'b1111;
	mem[3139] = 4'b1111;
	mem[3140] = 4'b1111;
	mem[3141] = 4'b1111;
	mem[3142] = 4'b1101;
	mem[3143] = 4'b0011;
	mem[3144] = 4'b0000;
	mem[3145] = 4'b0000;
	mem[3146] = 4'b0000;
	mem[3147] = 4'b0000;
	mem[3148] = 4'b0000;
	mem[3149] = 4'b0000;
	mem[3150] = 4'b0000;
	mem[3151] = 4'b0000;
	mem[3152] = 4'b0000;
	mem[3153] = 4'b0000;
	mem[3154] = 4'b0000;
	mem[3155] = 4'b0000;
	mem[3156] = 4'b0001;
	mem[3157] = 4'b0001;
	mem[3158] = 4'b0000;
	mem[3159] = 4'b0000;
	mem[3160] = 4'b0000;
	mem[3161] = 4'b0000;
	mem[3162] = 4'b0000;
	mem[3163] = 4'b0000;
	mem[3164] = 4'b0000;
	mem[3165] = 4'b0000;
	mem[3166] = 4'b0000;
	mem[3167] = 4'b0000;
	mem[3168] = 4'b0000;
	mem[3169] = 4'b0000;
	mem[3170] = 4'b0000;
	mem[3171] = 4'b0000;
	mem[3172] = 4'b0000;
	mem[3173] = 4'b0000;
	mem[3174] = 4'b0000;
	mem[3175] = 4'b0000;
	mem[3176] = 4'b0000;
	mem[3177] = 4'b0000;
	mem[3178] = 4'b0000;
	mem[3179] = 4'b0000;
	mem[3180] = 4'b0000;
	mem[3181] = 4'b0000;
	mem[3182] = 4'b0000;
	mem[3183] = 4'b0000;
	mem[3184] = 4'b0000;
	mem[3185] = 4'b0000;
	mem[3186] = 4'b0000;
	mem[3187] = 4'b0000;
	mem[3188] = 4'b0000;
	mem[3189] = 4'b0000;
	mem[3190] = 4'b0000;
	mem[3191] = 4'b0000;
	mem[3192] = 4'b0000;
	mem[3193] = 4'b0000;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b0111;
	mem[3204] = 4'b1100;
	mem[3205] = 4'b1101;
	mem[3206] = 4'b1110;
	mem[3207] = 4'b1110;
	mem[3208] = 4'b1110;
	mem[3209] = 4'b1110;
	mem[3210] = 4'b1110;
	mem[3211] = 4'b1110;
	mem[3212] = 4'b1110;
	mem[3213] = 4'b1110;
	mem[3214] = 4'b1110;
	mem[3215] = 4'b1110;
	mem[3216] = 4'b1101;
	mem[3217] = 4'b1100;
	mem[3218] = 4'b1100;
	mem[3219] = 4'b1110;
	mem[3220] = 4'b1111;
	mem[3221] = 4'b1111;
	mem[3222] = 4'b1111;
	mem[3223] = 4'b1111;
	mem[3224] = 4'b1101;
	mem[3225] = 4'b1110;
	mem[3226] = 4'b1111;
	mem[3227] = 4'b1111;
	mem[3228] = 4'b1111;
	mem[3229] = 4'b1111;
	mem[3230] = 4'b1111;
	mem[3231] = 4'b1111;
	mem[3232] = 4'b1111;
	mem[3233] = 4'b1111;
	mem[3234] = 4'b1111;
	mem[3235] = 4'b1111;
	mem[3236] = 4'b1111;
	mem[3237] = 4'b1111;
	mem[3238] = 4'b1111;
	mem[3239] = 4'b1111;
	mem[3240] = 4'b1111;
	mem[3241] = 4'b1111;
	mem[3242] = 4'b1111;
	mem[3243] = 4'b1111;
	mem[3244] = 4'b1111;
	mem[3245] = 4'b1111;
	mem[3246] = 4'b1111;
	mem[3247] = 4'b1111;
	mem[3248] = 4'b1111;
	mem[3249] = 4'b1111;
	mem[3250] = 4'b1111;
	mem[3251] = 4'b1111;
	mem[3252] = 4'b1111;
	mem[3253] = 4'b1111;
	mem[3254] = 4'b1111;
	mem[3255] = 4'b1111;
	mem[3256] = 4'b1111;
	mem[3257] = 4'b1111;
	mem[3258] = 4'b1111;
	mem[3259] = 4'b1111;
	mem[3260] = 4'b1111;
	mem[3261] = 4'b1111;
	mem[3262] = 4'b1111;
	mem[3263] = 4'b1111;
	mem[3264] = 4'b1111;
	mem[3265] = 4'b1111;
	mem[3266] = 4'b1111;
	mem[3267] = 4'b1111;
	mem[3268] = 4'b1111;
	mem[3269] = 4'b1111;
	mem[3270] = 4'b1111;
	mem[3271] = 4'b0011;
	mem[3272] = 4'b0000;
	mem[3273] = 4'b0000;
	mem[3274] = 4'b0000;
	mem[3275] = 4'b0000;
	mem[3276] = 4'b0001;
	mem[3277] = 4'b0000;
	mem[3278] = 4'b0000;
	mem[3279] = 4'b0000;
	mem[3280] = 4'b0000;
	mem[3281] = 4'b0000;
	mem[3282] = 4'b0000;
	mem[3283] = 4'b0001;
	mem[3284] = 4'b0001;
	mem[3285] = 4'b0000;
	mem[3286] = 4'b0000;
	mem[3287] = 4'b0000;
	mem[3288] = 4'b0000;
	mem[3289] = 4'b0000;
	mem[3290] = 4'b0000;
	mem[3291] = 4'b0000;
	mem[3292] = 4'b0000;
	mem[3293] = 4'b0000;
	mem[3294] = 4'b0000;
	mem[3295] = 4'b0000;
	mem[3296] = 4'b0000;
	mem[3297] = 4'b0000;
	mem[3298] = 4'b0000;
	mem[3299] = 4'b0000;
	mem[3300] = 4'b0000;
	mem[3301] = 4'b0000;
	mem[3302] = 4'b0000;
	mem[3303] = 4'b0000;
	mem[3304] = 4'b0000;
	mem[3305] = 4'b0000;
	mem[3306] = 4'b0000;
	mem[3307] = 4'b0000;
	mem[3308] = 4'b0000;
	mem[3309] = 4'b0000;
	mem[3310] = 4'b0000;
	mem[3311] = 4'b0000;
	mem[3312] = 4'b0000;
	mem[3313] = 4'b0000;
	mem[3314] = 4'b0000;
	mem[3315] = 4'b0000;
	mem[3316] = 4'b0000;
	mem[3317] = 4'b0000;
	mem[3318] = 4'b0000;
	mem[3319] = 4'b0000;
	mem[3320] = 4'b0000;
	mem[3321] = 4'b0000;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b0111;
	mem[3332] = 4'b1100;
	mem[3333] = 4'b1101;
	mem[3334] = 4'b1110;
	mem[3335] = 4'b1110;
	mem[3336] = 4'b1110;
	mem[3337] = 4'b1110;
	mem[3338] = 4'b1110;
	mem[3339] = 4'b1110;
	mem[3340] = 4'b1110;
	mem[3341] = 4'b1101;
	mem[3342] = 4'b1110;
	mem[3343] = 4'b1110;
	mem[3344] = 4'b1101;
	mem[3345] = 4'b1100;
	mem[3346] = 4'b1100;
	mem[3347] = 4'b1100;
	mem[3348] = 4'b1111;
	mem[3349] = 4'b1111;
	mem[3350] = 4'b1111;
	mem[3351] = 4'b1110;
	mem[3352] = 4'b1101;
	mem[3353] = 4'b1111;
	mem[3354] = 4'b1111;
	mem[3355] = 4'b1111;
	mem[3356] = 4'b1111;
	mem[3357] = 4'b1111;
	mem[3358] = 4'b1111;
	mem[3359] = 4'b1111;
	mem[3360] = 4'b1111;
	mem[3361] = 4'b1111;
	mem[3362] = 4'b1111;
	mem[3363] = 4'b1111;
	mem[3364] = 4'b1111;
	mem[3365] = 4'b1111;
	mem[3366] = 4'b1111;
	mem[3367] = 4'b1111;
	mem[3368] = 4'b1111;
	mem[3369] = 4'b1111;
	mem[3370] = 4'b1111;
	mem[3371] = 4'b1111;
	mem[3372] = 4'b1111;
	mem[3373] = 4'b1111;
	mem[3374] = 4'b1111;
	mem[3375] = 4'b1111;
	mem[3376] = 4'b1111;
	mem[3377] = 4'b1111;
	mem[3378] = 4'b1111;
	mem[3379] = 4'b1111;
	mem[3380] = 4'b1111;
	mem[3381] = 4'b1111;
	mem[3382] = 4'b1111;
	mem[3383] = 4'b1111;
	mem[3384] = 4'b1111;
	mem[3385] = 4'b1111;
	mem[3386] = 4'b1111;
	mem[3387] = 4'b1111;
	mem[3388] = 4'b1111;
	mem[3389] = 4'b1111;
	mem[3390] = 4'b1111;
	mem[3391] = 4'b1111;
	mem[3392] = 4'b1111;
	mem[3393] = 4'b1111;
	mem[3394] = 4'b1111;
	mem[3395] = 4'b1111;
	mem[3396] = 4'b1111;
	mem[3397] = 4'b1111;
	mem[3398] = 4'b1111;
	mem[3399] = 4'b0100;
	mem[3400] = 4'b0000;
	mem[3401] = 4'b0000;
	mem[3402] = 4'b0000;
	mem[3403] = 4'b0000;
	mem[3404] = 4'b0000;
	mem[3405] = 4'b0000;
	mem[3406] = 4'b0000;
	mem[3407] = 4'b0000;
	mem[3408] = 4'b0000;
	mem[3409] = 4'b0000;
	mem[3410] = 4'b0001;
	mem[3411] = 4'b0001;
	mem[3412] = 4'b0000;
	mem[3413] = 4'b0000;
	mem[3414] = 4'b0000;
	mem[3415] = 4'b0000;
	mem[3416] = 4'b0000;
	mem[3417] = 4'b0000;
	mem[3418] = 4'b0000;
	mem[3419] = 4'b0000;
	mem[3420] = 4'b0000;
	mem[3421] = 4'b0000;
	mem[3422] = 4'b0000;
	mem[3423] = 4'b0000;
	mem[3424] = 4'b0000;
	mem[3425] = 4'b0000;
	mem[3426] = 4'b0000;
	mem[3427] = 4'b0000;
	mem[3428] = 4'b0000;
	mem[3429] = 4'b0000;
	mem[3430] = 4'b0000;
	mem[3431] = 4'b0000;
	mem[3432] = 4'b0000;
	mem[3433] = 4'b0000;
	mem[3434] = 4'b0000;
	mem[3435] = 4'b0000;
	mem[3436] = 4'b0000;
	mem[3437] = 4'b0000;
	mem[3438] = 4'b0000;
	mem[3439] = 4'b0000;
	mem[3440] = 4'b0000;
	mem[3441] = 4'b0000;
	mem[3442] = 4'b0000;
	mem[3443] = 4'b0001;
	mem[3444] = 4'b0001;
	mem[3445] = 4'b0000;
	mem[3446] = 4'b0000;
	mem[3447] = 4'b0000;
	mem[3448] = 4'b0000;
	mem[3449] = 4'b0000;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b0111;
	mem[3460] = 4'b1100;
	mem[3461] = 4'b1101;
	mem[3462] = 4'b1110;
	mem[3463] = 4'b1110;
	mem[3464] = 4'b1110;
	mem[3465] = 4'b1110;
	mem[3466] = 4'b1110;
	mem[3467] = 4'b1101;
	mem[3468] = 4'b1100;
	mem[3469] = 4'b1100;
	mem[3470] = 4'b1100;
	mem[3471] = 4'b1101;
	mem[3472] = 4'b1110;
	mem[3473] = 4'b1101;
	mem[3474] = 4'b1100;
	mem[3475] = 4'b1100;
	mem[3476] = 4'b1101;
	mem[3477] = 4'b1110;
	mem[3478] = 4'b1110;
	mem[3479] = 4'b1101;
	mem[3480] = 4'b1110;
	mem[3481] = 4'b1111;
	mem[3482] = 4'b1111;
	mem[3483] = 4'b1111;
	mem[3484] = 4'b1111;
	mem[3485] = 4'b1111;
	mem[3486] = 4'b1111;
	mem[3487] = 4'b1111;
	mem[3488] = 4'b1111;
	mem[3489] = 4'b1111;
	mem[3490] = 4'b1111;
	mem[3491] = 4'b1111;
	mem[3492] = 4'b1111;
	mem[3493] = 4'b1111;
	mem[3494] = 4'b1111;
	mem[3495] = 4'b1111;
	mem[3496] = 4'b1111;
	mem[3497] = 4'b1111;
	mem[3498] = 4'b1111;
	mem[3499] = 4'b1111;
	mem[3500] = 4'b1111;
	mem[3501] = 4'b1111;
	mem[3502] = 4'b1111;
	mem[3503] = 4'b1111;
	mem[3504] = 4'b1111;
	mem[3505] = 4'b1111;
	mem[3506] = 4'b1111;
	mem[3507] = 4'b1111;
	mem[3508] = 4'b1111;
	mem[3509] = 4'b1111;
	mem[3510] = 4'b1111;
	mem[3511] = 4'b1111;
	mem[3512] = 4'b1111;
	mem[3513] = 4'b1111;
	mem[3514] = 4'b1111;
	mem[3515] = 4'b1111;
	mem[3516] = 4'b1111;
	mem[3517] = 4'b1111;
	mem[3518] = 4'b1111;
	mem[3519] = 4'b1111;
	mem[3520] = 4'b1111;
	mem[3521] = 4'b1111;
	mem[3522] = 4'b1111;
	mem[3523] = 4'b1111;
	mem[3524] = 4'b1101;
	mem[3525] = 4'b1111;
	mem[3526] = 4'b1111;
	mem[3527] = 4'b0100;
	mem[3528] = 4'b0000;
	mem[3529] = 4'b0000;
	mem[3530] = 4'b0000;
	mem[3531] = 4'b0000;
	mem[3532] = 4'b0000;
	mem[3533] = 4'b0000;
	mem[3534] = 4'b0000;
	mem[3535] = 4'b0000;
	mem[3536] = 4'b0000;
	mem[3537] = 4'b0001;
	mem[3538] = 4'b0001;
	mem[3539] = 4'b0000;
	mem[3540] = 4'b0000;
	mem[3541] = 4'b0000;
	mem[3542] = 4'b0000;
	mem[3543] = 4'b0000;
	mem[3544] = 4'b0000;
	mem[3545] = 4'b0000;
	mem[3546] = 4'b0000;
	mem[3547] = 4'b0000;
	mem[3548] = 4'b0000;
	mem[3549] = 4'b0000;
	mem[3550] = 4'b0000;
	mem[3551] = 4'b0000;
	mem[3552] = 4'b0000;
	mem[3553] = 4'b0000;
	mem[3554] = 4'b0000;
	mem[3555] = 4'b0000;
	mem[3556] = 4'b0000;
	mem[3557] = 4'b0000;
	mem[3558] = 4'b0000;
	mem[3559] = 4'b0000;
	mem[3560] = 4'b0000;
	mem[3561] = 4'b0000;
	mem[3562] = 4'b0000;
	mem[3563] = 4'b0000;
	mem[3564] = 4'b0000;
	mem[3565] = 4'b0000;
	mem[3566] = 4'b0000;
	mem[3567] = 4'b0000;
	mem[3568] = 4'b0000;
	mem[3569] = 4'b0000;
	mem[3570] = 4'b0001;
	mem[3571] = 4'b0001;
	mem[3572] = 4'b0000;
	mem[3573] = 4'b0000;
	mem[3574] = 4'b0000;
	mem[3575] = 4'b0000;
	mem[3576] = 4'b0000;
	mem[3577] = 4'b0000;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b0111;
	mem[3588] = 4'b1100;
	mem[3589] = 4'b1101;
	mem[3590] = 4'b1110;
	mem[3591] = 4'b1110;
	mem[3592] = 4'b1110;
	mem[3593] = 4'b1110;
	mem[3594] = 4'b1101;
	mem[3595] = 4'b1100;
	mem[3596] = 4'b1100;
	mem[3597] = 4'b1100;
	mem[3598] = 4'b1100;
	mem[3599] = 4'b1110;
	mem[3600] = 4'b1110;
	mem[3601] = 4'b1110;
	mem[3602] = 4'b1101;
	mem[3603] = 4'b1100;
	mem[3604] = 4'b1101;
	mem[3605] = 4'b1101;
	mem[3606] = 4'b1101;
	mem[3607] = 4'b1110;
	mem[3608] = 4'b1111;
	mem[3609] = 4'b1111;
	mem[3610] = 4'b1111;
	mem[3611] = 4'b1111;
	mem[3612] = 4'b1111;
	mem[3613] = 4'b1111;
	mem[3614] = 4'b1111;
	mem[3615] = 4'b1111;
	mem[3616] = 4'b1111;
	mem[3617] = 4'b1111;
	mem[3618] = 4'b1111;
	mem[3619] = 4'b1111;
	mem[3620] = 4'b1111;
	mem[3621] = 4'b1111;
	mem[3622] = 4'b1111;
	mem[3623] = 4'b1111;
	mem[3624] = 4'b1111;
	mem[3625] = 4'b1111;
	mem[3626] = 4'b1111;
	mem[3627] = 4'b1111;
	mem[3628] = 4'b1111;
	mem[3629] = 4'b1111;
	mem[3630] = 4'b1111;
	mem[3631] = 4'b1111;
	mem[3632] = 4'b1111;
	mem[3633] = 4'b1111;
	mem[3634] = 4'b1111;
	mem[3635] = 4'b1111;
	mem[3636] = 4'b1111;
	mem[3637] = 4'b1111;
	mem[3638] = 4'b1111;
	mem[3639] = 4'b1111;
	mem[3640] = 4'b1111;
	mem[3641] = 4'b1111;
	mem[3642] = 4'b1111;
	mem[3643] = 4'b1111;
	mem[3644] = 4'b1111;
	mem[3645] = 4'b1111;
	mem[3646] = 4'b1111;
	mem[3647] = 4'b1111;
	mem[3648] = 4'b1111;
	mem[3649] = 4'b1111;
	mem[3650] = 4'b1111;
	mem[3651] = 4'b1101;
	mem[3652] = 4'b1101;
	mem[3653] = 4'b1101;
	mem[3654] = 4'b1111;
	mem[3655] = 4'b0100;
	mem[3656] = 4'b0000;
	mem[3657] = 4'b0000;
	mem[3658] = 4'b0000;
	mem[3659] = 4'b0000;
	mem[3660] = 4'b0000;
	mem[3661] = 4'b0000;
	mem[3662] = 4'b0000;
	mem[3663] = 4'b0000;
	mem[3664] = 4'b0001;
	mem[3665] = 4'b0001;
	mem[3666] = 4'b0000;
	mem[3667] = 4'b0000;
	mem[3668] = 4'b0000;
	mem[3669] = 4'b0000;
	mem[3670] = 4'b0000;
	mem[3671] = 4'b0000;
	mem[3672] = 4'b0000;
	mem[3673] = 4'b0000;
	mem[3674] = 4'b0000;
	mem[3675] = 4'b0000;
	mem[3676] = 4'b0000;
	mem[3677] = 4'b0000;
	mem[3678] = 4'b0000;
	mem[3679] = 4'b0000;
	mem[3680] = 4'b0000;
	mem[3681] = 4'b0000;
	mem[3682] = 4'b0000;
	mem[3683] = 4'b0000;
	mem[3684] = 4'b0000;
	mem[3685] = 4'b0000;
	mem[3686] = 4'b0000;
	mem[3687] = 4'b0000;
	mem[3688] = 4'b0000;
	mem[3689] = 4'b0000;
	mem[3690] = 4'b0000;
	mem[3691] = 4'b0000;
	mem[3692] = 4'b0000;
	mem[3693] = 4'b0000;
	mem[3694] = 4'b0000;
	mem[3695] = 4'b0000;
	mem[3696] = 4'b0000;
	mem[3697] = 4'b0000;
	mem[3698] = 4'b0001;
	mem[3699] = 4'b0000;
	mem[3700] = 4'b0000;
	mem[3701] = 4'b0000;
	mem[3702] = 4'b0000;
	mem[3703] = 4'b0000;
	mem[3704] = 4'b0000;
	mem[3705] = 4'b0000;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b0111;
	mem[3716] = 4'b1100;
	mem[3717] = 4'b1101;
	mem[3718] = 4'b1110;
	mem[3719] = 4'b1110;
	mem[3720] = 4'b1110;
	mem[3721] = 4'b1101;
	mem[3722] = 4'b1100;
	mem[3723] = 4'b1100;
	mem[3724] = 4'b1101;
	mem[3725] = 4'b1110;
	mem[3726] = 4'b1110;
	mem[3727] = 4'b1110;
	mem[3728] = 4'b1110;
	mem[3729] = 4'b1101;
	mem[3730] = 4'b1110;
	mem[3731] = 4'b1110;
	mem[3732] = 4'b1111;
	mem[3733] = 4'b1111;
	mem[3734] = 4'b1111;
	mem[3735] = 4'b1111;
	mem[3736] = 4'b1111;
	mem[3737] = 4'b1111;
	mem[3738] = 4'b1111;
	mem[3739] = 4'b1111;
	mem[3740] = 4'b1111;
	mem[3741] = 4'b1111;
	mem[3742] = 4'b1111;
	mem[3743] = 4'b1111;
	mem[3744] = 4'b1111;
	mem[3745] = 4'b1111;
	mem[3746] = 4'b1111;
	mem[3747] = 4'b1111;
	mem[3748] = 4'b1111;
	mem[3749] = 4'b1111;
	mem[3750] = 4'b1111;
	mem[3751] = 4'b1111;
	mem[3752] = 4'b1111;
	mem[3753] = 4'b1111;
	mem[3754] = 4'b1111;
	mem[3755] = 4'b1111;
	mem[3756] = 4'b1111;
	mem[3757] = 4'b1111;
	mem[3758] = 4'b1111;
	mem[3759] = 4'b1111;
	mem[3760] = 4'b1111;
	mem[3761] = 4'b1111;
	mem[3762] = 4'b1111;
	mem[3763] = 4'b1111;
	mem[3764] = 4'b1111;
	mem[3765] = 4'b1111;
	mem[3766] = 4'b1111;
	mem[3767] = 4'b1111;
	mem[3768] = 4'b1111;
	mem[3769] = 4'b1111;
	mem[3770] = 4'b1111;
	mem[3771] = 4'b1111;
	mem[3772] = 4'b1111;
	mem[3773] = 4'b1111;
	mem[3774] = 4'b1111;
	mem[3775] = 4'b1111;
	mem[3776] = 4'b1111;
	mem[3777] = 4'b1111;
	mem[3778] = 4'b1101;
	mem[3779] = 4'b1101;
	mem[3780] = 4'b1101;
	mem[3781] = 4'b1101;
	mem[3782] = 4'b1110;
	mem[3783] = 4'b0100;
	mem[3784] = 4'b0000;
	mem[3785] = 4'b0000;
	mem[3786] = 4'b0000;
	mem[3787] = 4'b0000;
	mem[3788] = 4'b0000;
	mem[3789] = 4'b0000;
	mem[3790] = 4'b0000;
	mem[3791] = 4'b0001;
	mem[3792] = 4'b0001;
	mem[3793] = 4'b0000;
	mem[3794] = 4'b0000;
	mem[3795] = 4'b0000;
	mem[3796] = 4'b0000;
	mem[3797] = 4'b0000;
	mem[3798] = 4'b0000;
	mem[3799] = 4'b0000;
	mem[3800] = 4'b0000;
	mem[3801] = 4'b0000;
	mem[3802] = 4'b0000;
	mem[3803] = 4'b0000;
	mem[3804] = 4'b0000;
	mem[3805] = 4'b0000;
	mem[3806] = 4'b0000;
	mem[3807] = 4'b0000;
	mem[3808] = 4'b0000;
	mem[3809] = 4'b0000;
	mem[3810] = 4'b0000;
	mem[3811] = 4'b0000;
	mem[3812] = 4'b0000;
	mem[3813] = 4'b0000;
	mem[3814] = 4'b0000;
	mem[3815] = 4'b0000;
	mem[3816] = 4'b0000;
	mem[3817] = 4'b0000;
	mem[3818] = 4'b0000;
	mem[3819] = 4'b0000;
	mem[3820] = 4'b0000;
	mem[3821] = 4'b0000;
	mem[3822] = 4'b0000;
	mem[3823] = 4'b0000;
	mem[3824] = 4'b0000;
	mem[3825] = 4'b0000;
	mem[3826] = 4'b0000;
	mem[3827] = 4'b0000;
	mem[3828] = 4'b0000;
	mem[3829] = 4'b0000;
	mem[3830] = 4'b0000;
	mem[3831] = 4'b0000;
	mem[3832] = 4'b0000;
	mem[3833] = 4'b0000;
	mem[3834] = 4'b0001;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b0111;
	mem[3844] = 4'b1100;
	mem[3845] = 4'b1101;
	mem[3846] = 4'b1110;
	mem[3847] = 4'b1110;
	mem[3848] = 4'b1110;
	mem[3849] = 4'b1101;
	mem[3850] = 4'b1100;
	mem[3851] = 4'b1100;
	mem[3852] = 4'b1110;
	mem[3853] = 4'b1110;
	mem[3854] = 4'b1110;
	mem[3855] = 4'b1110;
	mem[3856] = 4'b1101;
	mem[3857] = 4'b1100;
	mem[3858] = 4'b1101;
	mem[3859] = 4'b1110;
	mem[3860] = 4'b1111;
	mem[3861] = 4'b1111;
	mem[3862] = 4'b1111;
	mem[3863] = 4'b1111;
	mem[3864] = 4'b1111;
	mem[3865] = 4'b1111;
	mem[3866] = 4'b1111;
	mem[3867] = 4'b1111;
	mem[3868] = 4'b1111;
	mem[3869] = 4'b1111;
	mem[3870] = 4'b1111;
	mem[3871] = 4'b1111;
	mem[3872] = 4'b1111;
	mem[3873] = 4'b1111;
	mem[3874] = 4'b1111;
	mem[3875] = 4'b1111;
	mem[3876] = 4'b1111;
	mem[3877] = 4'b1111;
	mem[3878] = 4'b1111;
	mem[3879] = 4'b1111;
	mem[3880] = 4'b1111;
	mem[3881] = 4'b1111;
	mem[3882] = 4'b1111;
	mem[3883] = 4'b1111;
	mem[3884] = 4'b1111;
	mem[3885] = 4'b1111;
	mem[3886] = 4'b1111;
	mem[3887] = 4'b1111;
	mem[3888] = 4'b1111;
	mem[3889] = 4'b1111;
	mem[3890] = 4'b1111;
	mem[3891] = 4'b1111;
	mem[3892] = 4'b1111;
	mem[3893] = 4'b1111;
	mem[3894] = 4'b1111;
	mem[3895] = 4'b1111;
	mem[3896] = 4'b1111;
	mem[3897] = 4'b1111;
	mem[3898] = 4'b1111;
	mem[3899] = 4'b1111;
	mem[3900] = 4'b1111;
	mem[3901] = 4'b1111;
	mem[3902] = 4'b1111;
	mem[3903] = 4'b1111;
	mem[3904] = 4'b1111;
	mem[3905] = 4'b1101;
	mem[3906] = 4'b1101;
	mem[3907] = 4'b1101;
	mem[3908] = 4'b1101;
	mem[3909] = 4'b1101;
	mem[3910] = 4'b1111;
	mem[3911] = 4'b0100;
	mem[3912] = 4'b0000;
	mem[3913] = 4'b0000;
	mem[3914] = 4'b0000;
	mem[3915] = 4'b0000;
	mem[3916] = 4'b0000;
	mem[3917] = 4'b0000;
	mem[3918] = 4'b0001;
	mem[3919] = 4'b0001;
	mem[3920] = 4'b0000;
	mem[3921] = 4'b0000;
	mem[3922] = 4'b0000;
	mem[3923] = 4'b0000;
	mem[3924] = 4'b0000;
	mem[3925] = 4'b0000;
	mem[3926] = 4'b0000;
	mem[3927] = 4'b0000;
	mem[3928] = 4'b0000;
	mem[3929] = 4'b0000;
	mem[3930] = 4'b0000;
	mem[3931] = 4'b0000;
	mem[3932] = 4'b0000;
	mem[3933] = 4'b0000;
	mem[3934] = 4'b0000;
	mem[3935] = 4'b0000;
	mem[3936] = 4'b0000;
	mem[3937] = 4'b0000;
	mem[3938] = 4'b0000;
	mem[3939] = 4'b0000;
	mem[3940] = 4'b0000;
	mem[3941] = 4'b0000;
	mem[3942] = 4'b0000;
	mem[3943] = 4'b0000;
	mem[3944] = 4'b0000;
	mem[3945] = 4'b0000;
	mem[3946] = 4'b0000;
	mem[3947] = 4'b0000;
	mem[3948] = 4'b0000;
	mem[3949] = 4'b0000;
	mem[3950] = 4'b0000;
	mem[3951] = 4'b0000;
	mem[3952] = 4'b0000;
	mem[3953] = 4'b0000;
	mem[3954] = 4'b0000;
	mem[3955] = 4'b0000;
	mem[3956] = 4'b0000;
	mem[3957] = 4'b0000;
	mem[3958] = 4'b0000;
	mem[3959] = 4'b0000;
	mem[3960] = 4'b0001;
	mem[3961] = 4'b0001;
	mem[3962] = 4'b0001;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b0111;
	mem[3972] = 4'b1011;
	mem[3973] = 4'b1100;
	mem[3974] = 4'b1110;
	mem[3975] = 4'b1110;
	mem[3976] = 4'b1110;
	mem[3977] = 4'b1101;
	mem[3978] = 4'b1100;
	mem[3979] = 4'b1100;
	mem[3980] = 4'b1110;
	mem[3981] = 4'b1110;
	mem[3982] = 4'b1110;
	mem[3983] = 4'b1110;
	mem[3984] = 4'b1101;
	mem[3985] = 4'b1100;
	mem[3986] = 4'b1100;
	mem[3987] = 4'b1110;
	mem[3988] = 4'b1111;
	mem[3989] = 4'b1111;
	mem[3990] = 4'b1111;
	mem[3991] = 4'b1111;
	mem[3992] = 4'b1111;
	mem[3993] = 4'b1111;
	mem[3994] = 4'b1111;
	mem[3995] = 4'b1111;
	mem[3996] = 4'b1111;
	mem[3997] = 4'b1111;
	mem[3998] = 4'b1111;
	mem[3999] = 4'b1111;
	mem[4000] = 4'b1111;
	mem[4001] = 4'b1111;
	mem[4002] = 4'b1111;
	mem[4003] = 4'b1111;
	mem[4004] = 4'b1111;
	mem[4005] = 4'b1111;
	mem[4006] = 4'b1111;
	mem[4007] = 4'b1111;
	mem[4008] = 4'b1111;
	mem[4009] = 4'b1111;
	mem[4010] = 4'b1111;
	mem[4011] = 4'b1111;
	mem[4012] = 4'b1111;
	mem[4013] = 4'b1111;
	mem[4014] = 4'b1111;
	mem[4015] = 4'b1111;
	mem[4016] = 4'b1111;
	mem[4017] = 4'b1111;
	mem[4018] = 4'b1111;
	mem[4019] = 4'b1111;
	mem[4020] = 4'b1111;
	mem[4021] = 4'b1111;
	mem[4022] = 4'b1111;
	mem[4023] = 4'b1111;
	mem[4024] = 4'b1111;
	mem[4025] = 4'b1111;
	mem[4026] = 4'b1111;
	mem[4027] = 4'b1111;
	mem[4028] = 4'b1111;
	mem[4029] = 4'b1111;
	mem[4030] = 4'b1111;
	mem[4031] = 4'b1110;
	mem[4032] = 4'b1101;
	mem[4033] = 4'b1101;
	mem[4034] = 4'b1101;
	mem[4035] = 4'b1101;
	mem[4036] = 4'b1101;
	mem[4037] = 4'b1111;
	mem[4038] = 4'b1111;
	mem[4039] = 4'b0100;
	mem[4040] = 4'b0000;
	mem[4041] = 4'b0000;
	mem[4042] = 4'b0000;
	mem[4043] = 4'b0000;
	mem[4044] = 4'b0000;
	mem[4045] = 4'b0001;
	mem[4046] = 4'b0001;
	mem[4047] = 4'b0000;
	mem[4048] = 4'b0000;
	mem[4049] = 4'b0000;
	mem[4050] = 4'b0000;
	mem[4051] = 4'b0000;
	mem[4052] = 4'b0000;
	mem[4053] = 4'b0000;
	mem[4054] = 4'b0000;
	mem[4055] = 4'b0000;
	mem[4056] = 4'b0000;
	mem[4057] = 4'b0000;
	mem[4058] = 4'b0000;
	mem[4059] = 4'b0000;
	mem[4060] = 4'b0000;
	mem[4061] = 4'b0000;
	mem[4062] = 4'b0000;
	mem[4063] = 4'b0000;
	mem[4064] = 4'b0000;
	mem[4065] = 4'b0000;
	mem[4066] = 4'b0000;
	mem[4067] = 4'b0000;
	mem[4068] = 4'b0000;
	mem[4069] = 4'b0000;
	mem[4070] = 4'b0000;
	mem[4071] = 4'b0000;
	mem[4072] = 4'b0000;
	mem[4073] = 4'b0000;
	mem[4074] = 4'b0000;
	mem[4075] = 4'b0000;
	mem[4076] = 4'b0000;
	mem[4077] = 4'b0000;
	mem[4078] = 4'b0000;
	mem[4079] = 4'b0000;
	mem[4080] = 4'b0000;
	mem[4081] = 4'b0000;
	mem[4082] = 4'b0000;
	mem[4083] = 4'b0000;
	mem[4084] = 4'b0000;
	mem[4085] = 4'b0000;
	mem[4086] = 4'b0000;
	mem[4087] = 4'b0000;
	mem[4088] = 4'b0001;
	mem[4089] = 4'b0000;
	mem[4090] = 4'b0000;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_2g (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0111;
	mem[4] = 4'b1011;
	mem[5] = 4'b1011;
	mem[6] = 4'b1101;
	mem[7] = 4'b1110;
	mem[8] = 4'b1110;
	mem[9] = 4'b1110;
	mem[10] = 4'b1100;
	mem[11] = 4'b1100;
	mem[12] = 4'b1101;
	mem[13] = 4'b1110;
	mem[14] = 4'b1110;
	mem[15] = 4'b1110;
	mem[16] = 4'b1101;
	mem[17] = 4'b1100;
	mem[18] = 4'b1100;
	mem[19] = 4'b1110;
	mem[20] = 4'b1111;
	mem[21] = 4'b1111;
	mem[22] = 4'b1111;
	mem[23] = 4'b1111;
	mem[24] = 4'b1111;
	mem[25] = 4'b1111;
	mem[26] = 4'b1111;
	mem[27] = 4'b1111;
	mem[28] = 4'b1111;
	mem[29] = 4'b1111;
	mem[30] = 4'b1111;
	mem[31] = 4'b1111;
	mem[32] = 4'b1111;
	mem[33] = 4'b1111;
	mem[34] = 4'b1111;
	mem[35] = 4'b1111;
	mem[36] = 4'b1111;
	mem[37] = 4'b1111;
	mem[38] = 4'b1111;
	mem[39] = 4'b1111;
	mem[40] = 4'b1111;
	mem[41] = 4'b1111;
	mem[42] = 4'b1111;
	mem[43] = 4'b1111;
	mem[44] = 4'b1111;
	mem[45] = 4'b1111;
	mem[46] = 4'b1111;
	mem[47] = 4'b1111;
	mem[48] = 4'b1111;
	mem[49] = 4'b1111;
	mem[50] = 4'b1111;
	mem[51] = 4'b1111;
	mem[52] = 4'b1111;
	mem[53] = 4'b1111;
	mem[54] = 4'b1111;
	mem[55] = 4'b1111;
	mem[56] = 4'b1111;
	mem[57] = 4'b1111;
	mem[58] = 4'b1111;
	mem[59] = 4'b1111;
	mem[60] = 4'b1111;
	mem[61] = 4'b1111;
	mem[62] = 4'b1111;
	mem[63] = 4'b1110;
	mem[64] = 4'b1101;
	mem[65] = 4'b1101;
	mem[66] = 4'b1101;
	mem[67] = 4'b1101;
	mem[68] = 4'b1111;
	mem[69] = 4'b1111;
	mem[70] = 4'b1111;
	mem[71] = 4'b0100;
	mem[72] = 4'b0000;
	mem[73] = 4'b0000;
	mem[74] = 4'b0000;
	mem[75] = 4'b0000;
	mem[76] = 4'b0000;
	mem[77] = 4'b0000;
	mem[78] = 4'b0000;
	mem[79] = 4'b0000;
	mem[80] = 4'b0000;
	mem[81] = 4'b0000;
	mem[82] = 4'b0000;
	mem[83] = 4'b0000;
	mem[84] = 4'b0000;
	mem[85] = 4'b0000;
	mem[86] = 4'b0000;
	mem[87] = 4'b0000;
	mem[88] = 4'b0000;
	mem[89] = 4'b0000;
	mem[90] = 4'b0000;
	mem[91] = 4'b0000;
	mem[92] = 4'b0000;
	mem[93] = 4'b0000;
	mem[94] = 4'b0000;
	mem[95] = 4'b0000;
	mem[96] = 4'b0000;
	mem[97] = 4'b0000;
	mem[98] = 4'b0000;
	mem[99] = 4'b0000;
	mem[100] = 4'b0000;
	mem[101] = 4'b0000;
	mem[102] = 4'b0000;
	mem[103] = 4'b0000;
	mem[104] = 4'b0000;
	mem[105] = 4'b0000;
	mem[106] = 4'b0000;
	mem[107] = 4'b0000;
	mem[108] = 4'b0000;
	mem[109] = 4'b0000;
	mem[110] = 4'b0000;
	mem[111] = 4'b0000;
	mem[112] = 4'b0000;
	mem[113] = 4'b0000;
	mem[114] = 4'b0000;
	mem[115] = 4'b0000;
	mem[116] = 4'b0000;
	mem[117] = 4'b0000;
	mem[118] = 4'b0000;
	mem[119] = 4'b0001;
	mem[120] = 4'b0001;
	mem[121] = 4'b0000;
	mem[122] = 4'b0000;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b1000;
	mem[132] = 4'b1100;
	mem[133] = 4'b1011;
	mem[134] = 4'b1100;
	mem[135] = 4'b1101;
	mem[136] = 4'b1110;
	mem[137] = 4'b1110;
	mem[138] = 4'b1101;
	mem[139] = 4'b1100;
	mem[140] = 4'b1100;
	mem[141] = 4'b1101;
	mem[142] = 4'b1101;
	mem[143] = 4'b1101;
	mem[144] = 4'b1100;
	mem[145] = 4'b1100;
	mem[146] = 4'b1101;
	mem[147] = 4'b1110;
	mem[148] = 4'b1111;
	mem[149] = 4'b1111;
	mem[150] = 4'b1111;
	mem[151] = 4'b1111;
	mem[152] = 4'b1111;
	mem[153] = 4'b1111;
	mem[154] = 4'b1111;
	mem[155] = 4'b1111;
	mem[156] = 4'b1111;
	mem[157] = 4'b1111;
	mem[158] = 4'b1111;
	mem[159] = 4'b1111;
	mem[160] = 4'b1111;
	mem[161] = 4'b1111;
	mem[162] = 4'b1111;
	mem[163] = 4'b1111;
	mem[164] = 4'b1111;
	mem[165] = 4'b1111;
	mem[166] = 4'b1111;
	mem[167] = 4'b1111;
	mem[168] = 4'b1111;
	mem[169] = 4'b1111;
	mem[170] = 4'b1111;
	mem[171] = 4'b1111;
	mem[172] = 4'b1111;
	mem[173] = 4'b1111;
	mem[174] = 4'b1111;
	mem[175] = 4'b1111;
	mem[176] = 4'b1111;
	mem[177] = 4'b1111;
	mem[178] = 4'b1111;
	mem[179] = 4'b1111;
	mem[180] = 4'b1111;
	mem[181] = 4'b1111;
	mem[182] = 4'b1110;
	mem[183] = 4'b1101;
	mem[184] = 4'b1101;
	mem[185] = 4'b1101;
	mem[186] = 4'b1110;
	mem[187] = 4'b1111;
	mem[188] = 4'b1111;
	mem[189] = 4'b1111;
	mem[190] = 4'b1111;
	mem[191] = 4'b1111;
	mem[192] = 4'b1110;
	mem[193] = 4'b1101;
	mem[194] = 4'b1101;
	mem[195] = 4'b1111;
	mem[196] = 4'b1111;
	mem[197] = 4'b1111;
	mem[198] = 4'b1111;
	mem[199] = 4'b0100;
	mem[200] = 4'b0000;
	mem[201] = 4'b0000;
	mem[202] = 4'b0000;
	mem[203] = 4'b0000;
	mem[204] = 4'b0000;
	mem[205] = 4'b0000;
	mem[206] = 4'b0000;
	mem[207] = 4'b0000;
	mem[208] = 4'b0000;
	mem[209] = 4'b0000;
	mem[210] = 4'b0000;
	mem[211] = 4'b0000;
	mem[212] = 4'b0000;
	mem[213] = 4'b0000;
	mem[214] = 4'b0000;
	mem[215] = 4'b0000;
	mem[216] = 4'b0000;
	mem[217] = 4'b0000;
	mem[218] = 4'b0000;
	mem[219] = 4'b0000;
	mem[220] = 4'b0000;
	mem[221] = 4'b0000;
	mem[222] = 4'b0000;
	mem[223] = 4'b0000;
	mem[224] = 4'b0000;
	mem[225] = 4'b0000;
	mem[226] = 4'b0000;
	mem[227] = 4'b0000;
	mem[228] = 4'b0000;
	mem[229] = 4'b0000;
	mem[230] = 4'b0000;
	mem[231] = 4'b0000;
	mem[232] = 4'b0000;
	mem[233] = 4'b0000;
	mem[234] = 4'b0000;
	mem[235] = 4'b0000;
	mem[236] = 4'b0000;
	mem[237] = 4'b0000;
	mem[238] = 4'b0000;
	mem[239] = 4'b0000;
	mem[240] = 4'b0000;
	mem[241] = 4'b0000;
	mem[242] = 4'b0000;
	mem[243] = 4'b0000;
	mem[244] = 4'b0001;
	mem[245] = 4'b0001;
	mem[246] = 4'b0001;
	mem[247] = 4'b0001;
	mem[248] = 4'b0000;
	mem[249] = 4'b0000;
	mem[250] = 4'b0000;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0111;
	mem[260] = 4'b1100;
	mem[261] = 4'b1100;
	mem[262] = 4'b1100;
	mem[263] = 4'b1100;
	mem[264] = 4'b1101;
	mem[265] = 4'b1110;
	mem[266] = 4'b1110;
	mem[267] = 4'b1101;
	mem[268] = 4'b1100;
	mem[269] = 4'b1100;
	mem[270] = 4'b1100;
	mem[271] = 4'b1100;
	mem[272] = 4'b1100;
	mem[273] = 4'b1101;
	mem[274] = 4'b1110;
	mem[275] = 4'b1110;
	mem[276] = 4'b1111;
	mem[277] = 4'b1111;
	mem[278] = 4'b1111;
	mem[279] = 4'b1111;
	mem[280] = 4'b1111;
	mem[281] = 4'b1111;
	mem[282] = 4'b1111;
	mem[283] = 4'b1111;
	mem[284] = 4'b1111;
	mem[285] = 4'b1111;
	mem[286] = 4'b1111;
	mem[287] = 4'b1111;
	mem[288] = 4'b1111;
	mem[289] = 4'b1111;
	mem[290] = 4'b1111;
	mem[291] = 4'b1111;
	mem[292] = 4'b1111;
	mem[293] = 4'b1111;
	mem[294] = 4'b1111;
	mem[295] = 4'b1111;
	mem[296] = 4'b1111;
	mem[297] = 4'b1111;
	mem[298] = 4'b1111;
	mem[299] = 4'b1111;
	mem[300] = 4'b1111;
	mem[301] = 4'b1111;
	mem[302] = 4'b1111;
	mem[303] = 4'b1111;
	mem[304] = 4'b1111;
	mem[305] = 4'b1111;
	mem[306] = 4'b1111;
	mem[307] = 4'b1111;
	mem[308] = 4'b1110;
	mem[309] = 4'b1101;
	mem[310] = 4'b1101;
	mem[311] = 4'b1101;
	mem[312] = 4'b1101;
	mem[313] = 4'b1101;
	mem[314] = 4'b1111;
	mem[315] = 4'b1111;
	mem[316] = 4'b1111;
	mem[317] = 4'b1111;
	mem[318] = 4'b1111;
	mem[319] = 4'b1111;
	mem[320] = 4'b1111;
	mem[321] = 4'b1110;
	mem[322] = 4'b1111;
	mem[323] = 4'b1111;
	mem[324] = 4'b1111;
	mem[325] = 4'b1111;
	mem[326] = 4'b1111;
	mem[327] = 4'b0100;
	mem[328] = 4'b0000;
	mem[329] = 4'b0000;
	mem[330] = 4'b0000;
	mem[331] = 4'b0000;
	mem[332] = 4'b0000;
	mem[333] = 4'b0000;
	mem[334] = 4'b0000;
	mem[335] = 4'b0000;
	mem[336] = 4'b0000;
	mem[337] = 4'b0000;
	mem[338] = 4'b0000;
	mem[339] = 4'b0000;
	mem[340] = 4'b0000;
	mem[341] = 4'b0000;
	mem[342] = 4'b0000;
	mem[343] = 4'b0000;
	mem[344] = 4'b0000;
	mem[345] = 4'b0000;
	mem[346] = 4'b0000;
	mem[347] = 4'b0000;
	mem[348] = 4'b0000;
	mem[349] = 4'b0000;
	mem[350] = 4'b0000;
	mem[351] = 4'b0000;
	mem[352] = 4'b0000;
	mem[353] = 4'b0000;
	mem[354] = 4'b0000;
	mem[355] = 4'b0000;
	mem[356] = 4'b0000;
	mem[357] = 4'b0000;
	mem[358] = 4'b0000;
	mem[359] = 4'b0000;
	mem[360] = 4'b0000;
	mem[361] = 4'b0000;
	mem[362] = 4'b0000;
	mem[363] = 4'b0001;
	mem[364] = 4'b0001;
	mem[365] = 4'b0000;
	mem[366] = 4'b0001;
	mem[367] = 4'b0000;
	mem[368] = 4'b0000;
	mem[369] = 4'b0000;
	mem[370] = 4'b0000;
	mem[371] = 4'b0000;
	mem[372] = 4'b0000;
	mem[373] = 4'b0000;
	mem[374] = 4'b0000;
	mem[375] = 4'b0000;
	mem[376] = 4'b0000;
	mem[377] = 4'b0000;
	mem[378] = 4'b0000;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0111;
	mem[388] = 4'b1100;
	mem[389] = 4'b1101;
	mem[390] = 4'b1101;
	mem[391] = 4'b1100;
	mem[392] = 4'b1100;
	mem[393] = 4'b1101;
	mem[394] = 4'b1110;
	mem[395] = 4'b1110;
	mem[396] = 4'b1101;
	mem[397] = 4'b1100;
	mem[398] = 4'b1100;
	mem[399] = 4'b1100;
	mem[400] = 4'b1101;
	mem[401] = 4'b1110;
	mem[402] = 4'b1110;
	mem[403] = 4'b1110;
	mem[404] = 4'b1111;
	mem[405] = 4'b1111;
	mem[406] = 4'b1111;
	mem[407] = 4'b1111;
	mem[408] = 4'b1111;
	mem[409] = 4'b1111;
	mem[410] = 4'b1111;
	mem[411] = 4'b1111;
	mem[412] = 4'b1111;
	mem[413] = 4'b1111;
	mem[414] = 4'b1111;
	mem[415] = 4'b1111;
	mem[416] = 4'b1111;
	mem[417] = 4'b1111;
	mem[418] = 4'b1111;
	mem[419] = 4'b1111;
	mem[420] = 4'b1111;
	mem[421] = 4'b1111;
	mem[422] = 4'b1111;
	mem[423] = 4'b1111;
	mem[424] = 4'b1111;
	mem[425] = 4'b1111;
	mem[426] = 4'b1111;
	mem[427] = 4'b1111;
	mem[428] = 4'b1111;
	mem[429] = 4'b1111;
	mem[430] = 4'b1111;
	mem[431] = 4'b1111;
	mem[432] = 4'b1111;
	mem[433] = 4'b1111;
	mem[434] = 4'b1111;
	mem[435] = 4'b1110;
	mem[436] = 4'b1101;
	mem[437] = 4'b1101;
	mem[438] = 4'b1101;
	mem[439] = 4'b1101;
	mem[440] = 4'b1101;
	mem[441] = 4'b1110;
	mem[442] = 4'b1111;
	mem[443] = 4'b1111;
	mem[444] = 4'b1111;
	mem[445] = 4'b1111;
	mem[446] = 4'b1111;
	mem[447] = 4'b1111;
	mem[448] = 4'b1111;
	mem[449] = 4'b1111;
	mem[450] = 4'b1111;
	mem[451] = 4'b1111;
	mem[452] = 4'b1111;
	mem[453] = 4'b1111;
	mem[454] = 4'b1111;
	mem[455] = 4'b0100;
	mem[456] = 4'b0000;
	mem[457] = 4'b0000;
	mem[458] = 4'b0000;
	mem[459] = 4'b0000;
	mem[460] = 4'b0000;
	mem[461] = 4'b0000;
	mem[462] = 4'b0000;
	mem[463] = 4'b0000;
	mem[464] = 4'b0000;
	mem[465] = 4'b0000;
	mem[466] = 4'b0000;
	mem[467] = 4'b0000;
	mem[468] = 4'b0000;
	mem[469] = 4'b0000;
	mem[470] = 4'b0000;
	mem[471] = 4'b0000;
	mem[472] = 4'b0000;
	mem[473] = 4'b0000;
	mem[474] = 4'b0000;
	mem[475] = 4'b0000;
	mem[476] = 4'b0000;
	mem[477] = 4'b0000;
	mem[478] = 4'b0000;
	mem[479] = 4'b0000;
	mem[480] = 4'b0000;
	mem[481] = 4'b0000;
	mem[482] = 4'b0000;
	mem[483] = 4'b0000;
	mem[484] = 4'b0000;
	mem[485] = 4'b0000;
	mem[486] = 4'b0000;
	mem[487] = 4'b0000;
	mem[488] = 4'b0000;
	mem[489] = 4'b0000;
	mem[490] = 4'b0000;
	mem[491] = 4'b0001;
	mem[492] = 4'b0000;
	mem[493] = 4'b0000;
	mem[494] = 4'b0000;
	mem[495] = 4'b0000;
	mem[496] = 4'b0000;
	mem[497] = 4'b0000;
	mem[498] = 4'b0000;
	mem[499] = 4'b0000;
	mem[500] = 4'b0000;
	mem[501] = 4'b0000;
	mem[502] = 4'b0000;
	mem[503] = 4'b0000;
	mem[504] = 4'b0000;
	mem[505] = 4'b0000;
	mem[506] = 4'b0000;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0111;
	mem[516] = 4'b1100;
	mem[517] = 4'b1101;
	mem[518] = 4'b1110;
	mem[519] = 4'b1101;
	mem[520] = 4'b1100;
	mem[521] = 4'b1100;
	mem[522] = 4'b1101;
	mem[523] = 4'b1110;
	mem[524] = 4'b1110;
	mem[525] = 4'b1110;
	mem[526] = 4'b1110;
	mem[527] = 4'b1110;
	mem[528] = 4'b1110;
	mem[529] = 4'b1110;
	mem[530] = 4'b1110;
	mem[531] = 4'b1101;
	mem[532] = 4'b1111;
	mem[533] = 4'b1111;
	mem[534] = 4'b1111;
	mem[535] = 4'b1111;
	mem[536] = 4'b1111;
	mem[537] = 4'b1111;
	mem[538] = 4'b1111;
	mem[539] = 4'b1111;
	mem[540] = 4'b1111;
	mem[541] = 4'b1111;
	mem[542] = 4'b1111;
	mem[543] = 4'b1111;
	mem[544] = 4'b1111;
	mem[545] = 4'b1111;
	mem[546] = 4'b1111;
	mem[547] = 4'b1111;
	mem[548] = 4'b1111;
	mem[549] = 4'b1111;
	mem[550] = 4'b1111;
	mem[551] = 4'b1111;
	mem[552] = 4'b1111;
	mem[553] = 4'b1111;
	mem[554] = 4'b1111;
	mem[555] = 4'b1111;
	mem[556] = 4'b1111;
	mem[557] = 4'b1111;
	mem[558] = 4'b1111;
	mem[559] = 4'b1111;
	mem[560] = 4'b1111;
	mem[561] = 4'b1111;
	mem[562] = 4'b1110;
	mem[563] = 4'b1101;
	mem[564] = 4'b1101;
	mem[565] = 4'b1101;
	mem[566] = 4'b1110;
	mem[567] = 4'b1111;
	mem[568] = 4'b1111;
	mem[569] = 4'b1111;
	mem[570] = 4'b1111;
	mem[571] = 4'b1111;
	mem[572] = 4'b1111;
	mem[573] = 4'b1110;
	mem[574] = 4'b1111;
	mem[575] = 4'b1111;
	mem[576] = 4'b1111;
	mem[577] = 4'b1111;
	mem[578] = 4'b1111;
	mem[579] = 4'b1111;
	mem[580] = 4'b1111;
	mem[581] = 4'b1111;
	mem[582] = 4'b1111;
	mem[583] = 4'b0100;
	mem[584] = 4'b0000;
	mem[585] = 4'b0000;
	mem[586] = 4'b0000;
	mem[587] = 4'b0000;
	mem[588] = 4'b0000;
	mem[589] = 4'b0000;
	mem[590] = 4'b0000;
	mem[591] = 4'b0000;
	mem[592] = 4'b0000;
	mem[593] = 4'b0000;
	mem[594] = 4'b0000;
	mem[595] = 4'b0000;
	mem[596] = 4'b0000;
	mem[597] = 4'b0000;
	mem[598] = 4'b0000;
	mem[599] = 4'b0000;
	mem[600] = 4'b0000;
	mem[601] = 4'b0000;
	mem[602] = 4'b0000;
	mem[603] = 4'b0000;
	mem[604] = 4'b0000;
	mem[605] = 4'b0000;
	mem[606] = 4'b0000;
	mem[607] = 4'b0000;
	mem[608] = 4'b0000;
	mem[609] = 4'b0000;
	mem[610] = 4'b0000;
	mem[611] = 4'b0000;
	mem[612] = 4'b0000;
	mem[613] = 4'b0000;
	mem[614] = 4'b0000;
	mem[615] = 4'b0000;
	mem[616] = 4'b0000;
	mem[617] = 4'b0000;
	mem[618] = 4'b0000;
	mem[619] = 4'b0000;
	mem[620] = 4'b0000;
	mem[621] = 4'b0000;
	mem[622] = 4'b0000;
	mem[623] = 4'b0000;
	mem[624] = 4'b0000;
	mem[625] = 4'b0000;
	mem[626] = 4'b0000;
	mem[627] = 4'b0001;
	mem[628] = 4'b0000;
	mem[629] = 4'b0000;
	mem[630] = 4'b0000;
	mem[631] = 4'b0000;
	mem[632] = 4'b0000;
	mem[633] = 4'b0000;
	mem[634] = 4'b0000;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0111;
	mem[644] = 4'b1100;
	mem[645] = 4'b1101;
	mem[646] = 4'b1110;
	mem[647] = 4'b1110;
	mem[648] = 4'b1101;
	mem[649] = 4'b1100;
	mem[650] = 4'b1100;
	mem[651] = 4'b1101;
	mem[652] = 4'b1110;
	mem[653] = 4'b1110;
	mem[654] = 4'b1110;
	mem[655] = 4'b1110;
	mem[656] = 4'b1110;
	mem[657] = 4'b1101;
	mem[658] = 4'b1100;
	mem[659] = 4'b1100;
	mem[660] = 4'b1111;
	mem[661] = 4'b1111;
	mem[662] = 4'b1111;
	mem[663] = 4'b1111;
	mem[664] = 4'b1111;
	mem[665] = 4'b1111;
	mem[666] = 4'b1111;
	mem[667] = 4'b1111;
	mem[668] = 4'b1111;
	mem[669] = 4'b1111;
	mem[670] = 4'b1111;
	mem[671] = 4'b1111;
	mem[672] = 4'b1111;
	mem[673] = 4'b1111;
	mem[674] = 4'b1111;
	mem[675] = 4'b1111;
	mem[676] = 4'b1111;
	mem[677] = 4'b1111;
	mem[678] = 4'b1111;
	mem[679] = 4'b1111;
	mem[680] = 4'b1111;
	mem[681] = 4'b1111;
	mem[682] = 4'b1111;
	mem[683] = 4'b1111;
	mem[684] = 4'b1111;
	mem[685] = 4'b1111;
	mem[686] = 4'b1111;
	mem[687] = 4'b1111;
	mem[688] = 4'b1111;
	mem[689] = 4'b1111;
	mem[690] = 4'b1101;
	mem[691] = 4'b1101;
	mem[692] = 4'b1101;
	mem[693] = 4'b1111;
	mem[694] = 4'b1111;
	mem[695] = 4'b1111;
	mem[696] = 4'b1111;
	mem[697] = 4'b1111;
	mem[698] = 4'b1110;
	mem[699] = 4'b1101;
	mem[700] = 4'b1101;
	mem[701] = 4'b1101;
	mem[702] = 4'b1101;
	mem[703] = 4'b1110;
	mem[704] = 4'b1111;
	mem[705] = 4'b1111;
	mem[706] = 4'b1111;
	mem[707] = 4'b1111;
	mem[708] = 4'b1111;
	mem[709] = 4'b1111;
	mem[710] = 4'b1111;
	mem[711] = 4'b0100;
	mem[712] = 4'b0000;
	mem[713] = 4'b0000;
	mem[714] = 4'b0000;
	mem[715] = 4'b0000;
	mem[716] = 4'b0000;
	mem[717] = 4'b0000;
	mem[718] = 4'b0000;
	mem[719] = 4'b0000;
	mem[720] = 4'b0000;
	mem[721] = 4'b0000;
	mem[722] = 4'b0000;
	mem[723] = 4'b0000;
	mem[724] = 4'b0000;
	mem[725] = 4'b0000;
	mem[726] = 4'b0000;
	mem[727] = 4'b0000;
	mem[728] = 4'b0000;
	mem[729] = 4'b0000;
	mem[730] = 4'b0000;
	mem[731] = 4'b0000;
	mem[732] = 4'b0000;
	mem[733] = 4'b0000;
	mem[734] = 4'b0000;
	mem[735] = 4'b0000;
	mem[736] = 4'b0000;
	mem[737] = 4'b0000;
	mem[738] = 4'b0000;
	mem[739] = 4'b0000;
	mem[740] = 4'b0000;
	mem[741] = 4'b0000;
	mem[742] = 4'b0000;
	mem[743] = 4'b0000;
	mem[744] = 4'b0000;
	mem[745] = 4'b0000;
	mem[746] = 4'b0000;
	mem[747] = 4'b0000;
	mem[748] = 4'b0000;
	mem[749] = 4'b0000;
	mem[750] = 4'b0000;
	mem[751] = 4'b0000;
	mem[752] = 4'b0000;
	mem[753] = 4'b0000;
	mem[754] = 4'b0001;
	mem[755] = 4'b0001;
	mem[756] = 4'b0000;
	mem[757] = 4'b0000;
	mem[758] = 4'b0000;
	mem[759] = 4'b0000;
	mem[760] = 4'b0000;
	mem[761] = 4'b0000;
	mem[762] = 4'b0000;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0111;
	mem[772] = 4'b1100;
	mem[773] = 4'b1101;
	mem[774] = 4'b1110;
	mem[775] = 4'b1110;
	mem[776] = 4'b1110;
	mem[777] = 4'b1101;
	mem[778] = 4'b1100;
	mem[779] = 4'b1100;
	mem[780] = 4'b1101;
	mem[781] = 4'b1110;
	mem[782] = 4'b1110;
	mem[783] = 4'b1110;
	mem[784] = 4'b1101;
	mem[785] = 4'b1100;
	mem[786] = 4'b1100;
	mem[787] = 4'b1100;
	mem[788] = 4'b1111;
	mem[789] = 4'b1111;
	mem[790] = 4'b1111;
	mem[791] = 4'b1111;
	mem[792] = 4'b1111;
	mem[793] = 4'b1111;
	mem[794] = 4'b1111;
	mem[795] = 4'b1111;
	mem[796] = 4'b1111;
	mem[797] = 4'b1111;
	mem[798] = 4'b1111;
	mem[799] = 4'b1111;
	mem[800] = 4'b1111;
	mem[801] = 4'b1111;
	mem[802] = 4'b1111;
	mem[803] = 4'b1111;
	mem[804] = 4'b1111;
	mem[805] = 4'b1111;
	mem[806] = 4'b1111;
	mem[807] = 4'b1111;
	mem[808] = 4'b1111;
	mem[809] = 4'b1111;
	mem[810] = 4'b1111;
	mem[811] = 4'b1111;
	mem[812] = 4'b1111;
	mem[813] = 4'b1111;
	mem[814] = 4'b1111;
	mem[815] = 4'b1111;
	mem[816] = 4'b1111;
	mem[817] = 4'b1110;
	mem[818] = 4'b1101;
	mem[819] = 4'b1101;
	mem[820] = 4'b1110;
	mem[821] = 4'b1111;
	mem[822] = 4'b1111;
	mem[823] = 4'b1111;
	mem[824] = 4'b1111;
	mem[825] = 4'b1101;
	mem[826] = 4'b1101;
	mem[827] = 4'b1101;
	mem[828] = 4'b1101;
	mem[829] = 4'b1101;
	mem[830] = 4'b1101;
	mem[831] = 4'b1101;
	mem[832] = 4'b1110;
	mem[833] = 4'b1111;
	mem[834] = 4'b1111;
	mem[835] = 4'b1111;
	mem[836] = 4'b1111;
	mem[837] = 4'b1111;
	mem[838] = 4'b1111;
	mem[839] = 4'b0100;
	mem[840] = 4'b0000;
	mem[841] = 4'b0000;
	mem[842] = 4'b0000;
	mem[843] = 4'b0000;
	mem[844] = 4'b0000;
	mem[845] = 4'b0000;
	mem[846] = 4'b0000;
	mem[847] = 4'b0000;
	mem[848] = 4'b0000;
	mem[849] = 4'b0000;
	mem[850] = 4'b0000;
	mem[851] = 4'b0000;
	mem[852] = 4'b0000;
	mem[853] = 4'b0000;
	mem[854] = 4'b0000;
	mem[855] = 4'b0000;
	mem[856] = 4'b0000;
	mem[857] = 4'b0000;
	mem[858] = 4'b0000;
	mem[859] = 4'b0000;
	mem[860] = 4'b0000;
	mem[861] = 4'b0000;
	mem[862] = 4'b0000;
	mem[863] = 4'b0000;
	mem[864] = 4'b0000;
	mem[865] = 4'b0000;
	mem[866] = 4'b0000;
	mem[867] = 4'b0000;
	mem[868] = 4'b0000;
	mem[869] = 4'b0000;
	mem[870] = 4'b0000;
	mem[871] = 4'b0000;
	mem[872] = 4'b0000;
	mem[873] = 4'b0000;
	mem[874] = 4'b0000;
	mem[875] = 4'b0000;
	mem[876] = 4'b0000;
	mem[877] = 4'b0000;
	mem[878] = 4'b0000;
	mem[879] = 4'b0000;
	mem[880] = 4'b0000;
	mem[881] = 4'b0000;
	mem[882] = 4'b0000;
	mem[883] = 4'b0000;
	mem[884] = 4'b0000;
	mem[885] = 4'b0000;
	mem[886] = 4'b0000;
	mem[887] = 4'b0000;
	mem[888] = 4'b0000;
	mem[889] = 4'b0000;
	mem[890] = 4'b0000;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0111;
	mem[900] = 4'b1100;
	mem[901] = 4'b1101;
	mem[902] = 4'b1110;
	mem[903] = 4'b1110;
	mem[904] = 4'b1110;
	mem[905] = 4'b1110;
	mem[906] = 4'b1101;
	mem[907] = 4'b1100;
	mem[908] = 4'b1101;
	mem[909] = 4'b1110;
	mem[910] = 4'b1101;
	mem[911] = 4'b1101;
	mem[912] = 4'b1100;
	mem[913] = 4'b1100;
	mem[914] = 4'b1100;
	mem[915] = 4'b1100;
	mem[916] = 4'b1111;
	mem[917] = 4'b1111;
	mem[918] = 4'b1111;
	mem[919] = 4'b1111;
	mem[920] = 4'b1111;
	mem[921] = 4'b1111;
	mem[922] = 4'b1111;
	mem[923] = 4'b1111;
	mem[924] = 4'b1111;
	mem[925] = 4'b1111;
	mem[926] = 4'b1111;
	mem[927] = 4'b1111;
	mem[928] = 4'b1111;
	mem[929] = 4'b1111;
	mem[930] = 4'b1111;
	mem[931] = 4'b1111;
	mem[932] = 4'b1111;
	mem[933] = 4'b1111;
	mem[934] = 4'b1111;
	mem[935] = 4'b1111;
	mem[936] = 4'b1111;
	mem[937] = 4'b1111;
	mem[938] = 4'b1111;
	mem[939] = 4'b1111;
	mem[940] = 4'b1111;
	mem[941] = 4'b1111;
	mem[942] = 4'b1111;
	mem[943] = 4'b1111;
	mem[944] = 4'b1111;
	mem[945] = 4'b1110;
	mem[946] = 4'b1101;
	mem[947] = 4'b1101;
	mem[948] = 4'b1111;
	mem[949] = 4'b1111;
	mem[950] = 4'b1111;
	mem[951] = 4'b1110;
	mem[952] = 4'b1101;
	mem[953] = 4'b1101;
	mem[954] = 4'b1101;
	mem[955] = 4'b1101;
	mem[956] = 4'b1101;
	mem[957] = 4'b1101;
	mem[958] = 4'b1101;
	mem[959] = 4'b1101;
	mem[960] = 4'b1101;
	mem[961] = 4'b1111;
	mem[962] = 4'b1111;
	mem[963] = 4'b1111;
	mem[964] = 4'b1111;
	mem[965] = 4'b1111;
	mem[966] = 4'b1111;
	mem[967] = 4'b0100;
	mem[968] = 4'b0000;
	mem[969] = 4'b0000;
	mem[970] = 4'b0000;
	mem[971] = 4'b0000;
	mem[972] = 4'b0000;
	mem[973] = 4'b0000;
	mem[974] = 4'b0000;
	mem[975] = 4'b0000;
	mem[976] = 4'b0000;
	mem[977] = 4'b0000;
	mem[978] = 4'b0000;
	mem[979] = 4'b0000;
	mem[980] = 4'b0000;
	mem[981] = 4'b0000;
	mem[982] = 4'b0000;
	mem[983] = 4'b0000;
	mem[984] = 4'b0000;
	mem[985] = 4'b0000;
	mem[986] = 4'b0000;
	mem[987] = 4'b0000;
	mem[988] = 4'b0000;
	mem[989] = 4'b0000;
	mem[990] = 4'b0000;
	mem[991] = 4'b0000;
	mem[992] = 4'b0000;
	mem[993] = 4'b0000;
	mem[994] = 4'b0000;
	mem[995] = 4'b0000;
	mem[996] = 4'b0000;
	mem[997] = 4'b0000;
	mem[998] = 4'b0000;
	mem[999] = 4'b0000;
	mem[1000] = 4'b0000;
	mem[1001] = 4'b0000;
	mem[1002] = 4'b0000;
	mem[1003] = 4'b0000;
	mem[1004] = 4'b0000;
	mem[1005] = 4'b0000;
	mem[1006] = 4'b0000;
	mem[1007] = 4'b0000;
	mem[1008] = 4'b0000;
	mem[1009] = 4'b0000;
	mem[1010] = 4'b0000;
	mem[1011] = 4'b0000;
	mem[1012] = 4'b0000;
	mem[1013] = 4'b0000;
	mem[1014] = 4'b0000;
	mem[1015] = 4'b0000;
	mem[1016] = 4'b0000;
	mem[1017] = 4'b0000;
	mem[1018] = 4'b0000;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0111;
	mem[1028] = 4'b1100;
	mem[1029] = 4'b1101;
	mem[1030] = 4'b1110;
	mem[1031] = 4'b1110;
	mem[1032] = 4'b1110;
	mem[1033] = 4'b1110;
	mem[1034] = 4'b1110;
	mem[1035] = 4'b1101;
	mem[1036] = 4'b1110;
	mem[1037] = 4'b1101;
	mem[1038] = 4'b1100;
	mem[1039] = 4'b1100;
	mem[1040] = 4'b1100;
	mem[1041] = 4'b1100;
	mem[1042] = 4'b1100;
	mem[1043] = 4'b1100;
	mem[1044] = 4'b1111;
	mem[1045] = 4'b1111;
	mem[1046] = 4'b1111;
	mem[1047] = 4'b1111;
	mem[1048] = 4'b1111;
	mem[1049] = 4'b1111;
	mem[1050] = 4'b1111;
	mem[1051] = 4'b1111;
	mem[1052] = 4'b1111;
	mem[1053] = 4'b1111;
	mem[1054] = 4'b1111;
	mem[1055] = 4'b1111;
	mem[1056] = 4'b1111;
	mem[1057] = 4'b1111;
	mem[1058] = 4'b1111;
	mem[1059] = 4'b1111;
	mem[1060] = 4'b1111;
	mem[1061] = 4'b1111;
	mem[1062] = 4'b1111;
	mem[1063] = 4'b1111;
	mem[1064] = 4'b1111;
	mem[1065] = 4'b1111;
	mem[1066] = 4'b1111;
	mem[1067] = 4'b1111;
	mem[1068] = 4'b1111;
	mem[1069] = 4'b1111;
	mem[1070] = 4'b1111;
	mem[1071] = 4'b1111;
	mem[1072] = 4'b1111;
	mem[1073] = 4'b1110;
	mem[1074] = 4'b1101;
	mem[1075] = 4'b1101;
	mem[1076] = 4'b1110;
	mem[1077] = 4'b1110;
	mem[1078] = 4'b1101;
	mem[1079] = 4'b1101;
	mem[1080] = 4'b1101;
	mem[1081] = 4'b1101;
	mem[1082] = 4'b1101;
	mem[1083] = 4'b1101;
	mem[1084] = 4'b1110;
	mem[1085] = 4'b1110;
	mem[1086] = 4'b1101;
	mem[1087] = 4'b1101;
	mem[1088] = 4'b1101;
	mem[1089] = 4'b1111;
	mem[1090] = 4'b1111;
	mem[1091] = 4'b1111;
	mem[1092] = 4'b1111;
	mem[1093] = 4'b1111;
	mem[1094] = 4'b1111;
	mem[1095] = 4'b0100;
	mem[1096] = 4'b0000;
	mem[1097] = 4'b0000;
	mem[1098] = 4'b0000;
	mem[1099] = 4'b0000;
	mem[1100] = 4'b0000;
	mem[1101] = 4'b0000;
	mem[1102] = 4'b0000;
	mem[1103] = 4'b0000;
	mem[1104] = 4'b0000;
	mem[1105] = 4'b0000;
	mem[1106] = 4'b0000;
	mem[1107] = 4'b0000;
	mem[1108] = 4'b0000;
	mem[1109] = 4'b0000;
	mem[1110] = 4'b0000;
	mem[1111] = 4'b0000;
	mem[1112] = 4'b0000;
	mem[1113] = 4'b0000;
	mem[1114] = 4'b0000;
	mem[1115] = 4'b0000;
	mem[1116] = 4'b0000;
	mem[1117] = 4'b0000;
	mem[1118] = 4'b0000;
	mem[1119] = 4'b0000;
	mem[1120] = 4'b0000;
	mem[1121] = 4'b0000;
	mem[1122] = 4'b0000;
	mem[1123] = 4'b0000;
	mem[1124] = 4'b0000;
	mem[1125] = 4'b0001;
	mem[1126] = 4'b0000;
	mem[1127] = 4'b0000;
	mem[1128] = 4'b0000;
	mem[1129] = 4'b0000;
	mem[1130] = 4'b0000;
	mem[1131] = 4'b0000;
	mem[1132] = 4'b0000;
	mem[1133] = 4'b0000;
	mem[1134] = 4'b0000;
	mem[1135] = 4'b0001;
	mem[1136] = 4'b0000;
	mem[1137] = 4'b0000;
	mem[1138] = 4'b0000;
	mem[1139] = 4'b0000;
	mem[1140] = 4'b0000;
	mem[1141] = 4'b0000;
	mem[1142] = 4'b0000;
	mem[1143] = 4'b0000;
	mem[1144] = 4'b0000;
	mem[1145] = 4'b0000;
	mem[1146] = 4'b0000;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0111;
	mem[1156] = 4'b1100;
	mem[1157] = 4'b1101;
	mem[1158] = 4'b1110;
	mem[1159] = 4'b1110;
	mem[1160] = 4'b1110;
	mem[1161] = 4'b1110;
	mem[1162] = 4'b1110;
	mem[1163] = 4'b1110;
	mem[1164] = 4'b1101;
	mem[1165] = 4'b1100;
	mem[1166] = 4'b1100;
	mem[1167] = 4'b1100;
	mem[1168] = 4'b1100;
	mem[1169] = 4'b1100;
	mem[1170] = 4'b1100;
	mem[1171] = 4'b1100;
	mem[1172] = 4'b1111;
	mem[1173] = 4'b1111;
	mem[1174] = 4'b1111;
	mem[1175] = 4'b1111;
	mem[1176] = 4'b1111;
	mem[1177] = 4'b1111;
	mem[1178] = 4'b1111;
	mem[1179] = 4'b1111;
	mem[1180] = 4'b1111;
	mem[1181] = 4'b1111;
	mem[1182] = 4'b1111;
	mem[1183] = 4'b1111;
	mem[1184] = 4'b1111;
	mem[1185] = 4'b1111;
	mem[1186] = 4'b1111;
	mem[1187] = 4'b1111;
	mem[1188] = 4'b1111;
	mem[1189] = 4'b1111;
	mem[1190] = 4'b1111;
	mem[1191] = 4'b1111;
	mem[1192] = 4'b1111;
	mem[1193] = 4'b1111;
	mem[1194] = 4'b1111;
	mem[1195] = 4'b1111;
	mem[1196] = 4'b1111;
	mem[1197] = 4'b1111;
	mem[1198] = 4'b1111;
	mem[1199] = 4'b1111;
	mem[1200] = 4'b1111;
	mem[1201] = 4'b1110;
	mem[1202] = 4'b1101;
	mem[1203] = 4'b1101;
	mem[1204] = 4'b1101;
	mem[1205] = 4'b1101;
	mem[1206] = 4'b1101;
	mem[1207] = 4'b1101;
	mem[1208] = 4'b1101;
	mem[1209] = 4'b1101;
	mem[1210] = 4'b1110;
	mem[1211] = 4'b1111;
	mem[1212] = 4'b1111;
	mem[1213] = 4'b1111;
	mem[1214] = 4'b1110;
	mem[1215] = 4'b1101;
	mem[1216] = 4'b1101;
	mem[1217] = 4'b1111;
	mem[1218] = 4'b1111;
	mem[1219] = 4'b1111;
	mem[1220] = 4'b1111;
	mem[1221] = 4'b1111;
	mem[1222] = 4'b1111;
	mem[1223] = 4'b0100;
	mem[1224] = 4'b0000;
	mem[1225] = 4'b0000;
	mem[1226] = 4'b0000;
	mem[1227] = 4'b0000;
	mem[1228] = 4'b0000;
	mem[1229] = 4'b0000;
	mem[1230] = 4'b0000;
	mem[1231] = 4'b0000;
	mem[1232] = 4'b0000;
	mem[1233] = 4'b0000;
	mem[1234] = 4'b0000;
	mem[1235] = 4'b0000;
	mem[1236] = 4'b0000;
	mem[1237] = 4'b0000;
	mem[1238] = 4'b0000;
	mem[1239] = 4'b0000;
	mem[1240] = 4'b0000;
	mem[1241] = 4'b0000;
	mem[1242] = 4'b0000;
	mem[1243] = 4'b0000;
	mem[1244] = 4'b0000;
	mem[1245] = 4'b0000;
	mem[1246] = 4'b0000;
	mem[1247] = 4'b0000;
	mem[1248] = 4'b0000;
	mem[1249] = 4'b0000;
	mem[1250] = 4'b0000;
	mem[1251] = 4'b0000;
	mem[1252] = 4'b0001;
	mem[1253] = 4'b0001;
	mem[1254] = 4'b0000;
	mem[1255] = 4'b0000;
	mem[1256] = 4'b0000;
	mem[1257] = 4'b0000;
	mem[1258] = 4'b0000;
	mem[1259] = 4'b0000;
	mem[1260] = 4'b0000;
	mem[1261] = 4'b0000;
	mem[1262] = 4'b0001;
	mem[1263] = 4'b0001;
	mem[1264] = 4'b0000;
	mem[1265] = 4'b0000;
	mem[1266] = 4'b0000;
	mem[1267] = 4'b0000;
	mem[1268] = 4'b0000;
	mem[1269] = 4'b0000;
	mem[1270] = 4'b0000;
	mem[1271] = 4'b0000;
	mem[1272] = 4'b0000;
	mem[1273] = 4'b0000;
	mem[1274] = 4'b0000;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0111;
	mem[1284] = 4'b1100;
	mem[1285] = 4'b1101;
	mem[1286] = 4'b1110;
	mem[1287] = 4'b1110;
	mem[1288] = 4'b1110;
	mem[1289] = 4'b1110;
	mem[1290] = 4'b1110;
	mem[1291] = 4'b1101;
	mem[1292] = 4'b1100;
	mem[1293] = 4'b1100;
	mem[1294] = 4'b1100;
	mem[1295] = 4'b1100;
	mem[1296] = 4'b1100;
	mem[1297] = 4'b1100;
	mem[1298] = 4'b1100;
	mem[1299] = 4'b1100;
	mem[1300] = 4'b1111;
	mem[1301] = 4'b1111;
	mem[1302] = 4'b1111;
	mem[1303] = 4'b1111;
	mem[1304] = 4'b1111;
	mem[1305] = 4'b1111;
	mem[1306] = 4'b1111;
	mem[1307] = 4'b1111;
	mem[1308] = 4'b1111;
	mem[1309] = 4'b1111;
	mem[1310] = 4'b1111;
	mem[1311] = 4'b1111;
	mem[1312] = 4'b1111;
	mem[1313] = 4'b1111;
	mem[1314] = 4'b1111;
	mem[1315] = 4'b1111;
	mem[1316] = 4'b1111;
	mem[1317] = 4'b1111;
	mem[1318] = 4'b1111;
	mem[1319] = 4'b1111;
	mem[1320] = 4'b1111;
	mem[1321] = 4'b1111;
	mem[1322] = 4'b1111;
	mem[1323] = 4'b1111;
	mem[1324] = 4'b1111;
	mem[1325] = 4'b1111;
	mem[1326] = 4'b1111;
	mem[1327] = 4'b1111;
	mem[1328] = 4'b1111;
	mem[1329] = 4'b1111;
	mem[1330] = 4'b1101;
	mem[1331] = 4'b1101;
	mem[1332] = 4'b1101;
	mem[1333] = 4'b1101;
	mem[1334] = 4'b1101;
	mem[1335] = 4'b1101;
	mem[1336] = 4'b1101;
	mem[1337] = 4'b1110;
	mem[1338] = 4'b1111;
	mem[1339] = 4'b1111;
	mem[1340] = 4'b1111;
	mem[1341] = 4'b1111;
	mem[1342] = 4'b1110;
	mem[1343] = 4'b1101;
	mem[1344] = 4'b1101;
	mem[1345] = 4'b1111;
	mem[1346] = 4'b1111;
	mem[1347] = 4'b1111;
	mem[1348] = 4'b1111;
	mem[1349] = 4'b1111;
	mem[1350] = 4'b1111;
	mem[1351] = 4'b0100;
	mem[1352] = 4'b0000;
	mem[1353] = 4'b0000;
	mem[1354] = 4'b0000;
	mem[1355] = 4'b0000;
	mem[1356] = 4'b0000;
	mem[1357] = 4'b0000;
	mem[1358] = 4'b0000;
	mem[1359] = 4'b0000;
	mem[1360] = 4'b0000;
	mem[1361] = 4'b0000;
	mem[1362] = 4'b0000;
	mem[1363] = 4'b0000;
	mem[1364] = 4'b0000;
	mem[1365] = 4'b0000;
	mem[1366] = 4'b0000;
	mem[1367] = 4'b0000;
	mem[1368] = 4'b0000;
	mem[1369] = 4'b0000;
	mem[1370] = 4'b0000;
	mem[1371] = 4'b0000;
	mem[1372] = 4'b0000;
	mem[1373] = 4'b0000;
	mem[1374] = 4'b0000;
	mem[1375] = 4'b0000;
	mem[1376] = 4'b0000;
	mem[1377] = 4'b0000;
	mem[1378] = 4'b0000;
	mem[1379] = 4'b0000;
	mem[1380] = 4'b0001;
	mem[1381] = 4'b0000;
	mem[1382] = 4'b0000;
	mem[1383] = 4'b0000;
	mem[1384] = 4'b0001;
	mem[1385] = 4'b0000;
	mem[1386] = 4'b0000;
	mem[1387] = 4'b0000;
	mem[1388] = 4'b0000;
	mem[1389] = 4'b0000;
	mem[1390] = 4'b0000;
	mem[1391] = 4'b0000;
	mem[1392] = 4'b0000;
	mem[1393] = 4'b0000;
	mem[1394] = 4'b0000;
	mem[1395] = 4'b0000;
	mem[1396] = 4'b0000;
	mem[1397] = 4'b0000;
	mem[1398] = 4'b0000;
	mem[1399] = 4'b0000;
	mem[1400] = 4'b0000;
	mem[1401] = 4'b0000;
	mem[1402] = 4'b0000;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0111;
	mem[1412] = 4'b1100;
	mem[1413] = 4'b1101;
	mem[1414] = 4'b1110;
	mem[1415] = 4'b1110;
	mem[1416] = 4'b1110;
	mem[1417] = 4'b1101;
	mem[1418] = 4'b1100;
	mem[1419] = 4'b1100;
	mem[1420] = 4'b1100;
	mem[1421] = 4'b1100;
	mem[1422] = 4'b1100;
	mem[1423] = 4'b1100;
	mem[1424] = 4'b1100;
	mem[1425] = 4'b1100;
	mem[1426] = 4'b1100;
	mem[1427] = 4'b1100;
	mem[1428] = 4'b1111;
	mem[1429] = 4'b1111;
	mem[1430] = 4'b1111;
	mem[1431] = 4'b1111;
	mem[1432] = 4'b1111;
	mem[1433] = 4'b1111;
	mem[1434] = 4'b1111;
	mem[1435] = 4'b1111;
	mem[1436] = 4'b1111;
	mem[1437] = 4'b1111;
	mem[1438] = 4'b1111;
	mem[1439] = 4'b1111;
	mem[1440] = 4'b1111;
	mem[1441] = 4'b1111;
	mem[1442] = 4'b1111;
	mem[1443] = 4'b1111;
	mem[1444] = 4'b1111;
	mem[1445] = 4'b1111;
	mem[1446] = 4'b1111;
	mem[1447] = 4'b1111;
	mem[1448] = 4'b1111;
	mem[1449] = 4'b1111;
	mem[1450] = 4'b1111;
	mem[1451] = 4'b1111;
	mem[1452] = 4'b1111;
	mem[1453] = 4'b1111;
	mem[1454] = 4'b1111;
	mem[1455] = 4'b1111;
	mem[1456] = 4'b1111;
	mem[1457] = 4'b1111;
	mem[1458] = 4'b1111;
	mem[1459] = 4'b1110;
	mem[1460] = 4'b1101;
	mem[1461] = 4'b1101;
	mem[1462] = 4'b1110;
	mem[1463] = 4'b1110;
	mem[1464] = 4'b1111;
	mem[1465] = 4'b1111;
	mem[1466] = 4'b1111;
	mem[1467] = 4'b1111;
	mem[1468] = 4'b1111;
	mem[1469] = 4'b1110;
	mem[1470] = 4'b1101;
	mem[1471] = 4'b1101;
	mem[1472] = 4'b1110;
	mem[1473] = 4'b1111;
	mem[1474] = 4'b1111;
	mem[1475] = 4'b1111;
	mem[1476] = 4'b1111;
	mem[1477] = 4'b1111;
	mem[1478] = 4'b1111;
	mem[1479] = 4'b0100;
	mem[1480] = 4'b0000;
	mem[1481] = 4'b0000;
	mem[1482] = 4'b0000;
	mem[1483] = 4'b0000;
	mem[1484] = 4'b0000;
	mem[1485] = 4'b0000;
	mem[1486] = 4'b0000;
	mem[1487] = 4'b0000;
	mem[1488] = 4'b0000;
	mem[1489] = 4'b0000;
	mem[1490] = 4'b0000;
	mem[1491] = 4'b0000;
	mem[1492] = 4'b0000;
	mem[1493] = 4'b0000;
	mem[1494] = 4'b0000;
	mem[1495] = 4'b0000;
	mem[1496] = 4'b0000;
	mem[1497] = 4'b0000;
	mem[1498] = 4'b0000;
	mem[1499] = 4'b0000;
	mem[1500] = 4'b0000;
	mem[1501] = 4'b0000;
	mem[1502] = 4'b0000;
	mem[1503] = 4'b0000;
	mem[1504] = 4'b0000;
	mem[1505] = 4'b0000;
	mem[1506] = 4'b0000;
	mem[1507] = 4'b0000;
	mem[1508] = 4'b0001;
	mem[1509] = 4'b0000;
	mem[1510] = 4'b0000;
	mem[1511] = 4'b0001;
	mem[1512] = 4'b0001;
	mem[1513] = 4'b0000;
	mem[1514] = 4'b0000;
	mem[1515] = 4'b0000;
	mem[1516] = 4'b0001;
	mem[1517] = 4'b0000;
	mem[1518] = 4'b0000;
	mem[1519] = 4'b0000;
	mem[1520] = 4'b0000;
	mem[1521] = 4'b0000;
	mem[1522] = 4'b0000;
	mem[1523] = 4'b0000;
	mem[1524] = 4'b0000;
	mem[1525] = 4'b0000;
	mem[1526] = 4'b0000;
	mem[1527] = 4'b0000;
	mem[1528] = 4'b0000;
	mem[1529] = 4'b0000;
	mem[1530] = 4'b0000;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0001;
	mem[1540] = 4'b0001;
	mem[1541] = 4'b0101;
	mem[1542] = 4'b1000;
	mem[1543] = 4'b1000;
	mem[1544] = 4'b0101;
	mem[1545] = 4'b0001;
	mem[1546] = 4'b0001;
	mem[1547] = 4'b0001;
	mem[1548] = 4'b0001;
	mem[1549] = 4'b0001;
	mem[1550] = 4'b0001;
	mem[1551] = 4'b0001;
	mem[1552] = 4'b0001;
	mem[1553] = 4'b0001;
	mem[1554] = 4'b0001;
	mem[1555] = 4'b0001;
	mem[1556] = 4'b0001;
	mem[1557] = 4'b0010;
	mem[1558] = 4'b0010;
	mem[1559] = 4'b0010;
	mem[1560] = 4'b0010;
	mem[1561] = 4'b0010;
	mem[1562] = 4'b0010;
	mem[1563] = 4'b0010;
	mem[1564] = 4'b0010;
	mem[1565] = 4'b0010;
	mem[1566] = 4'b0010;
	mem[1567] = 4'b0010;
	mem[1568] = 4'b0010;
	mem[1569] = 4'b0010;
	mem[1570] = 4'b0010;
	mem[1571] = 4'b0010;
	mem[1572] = 4'b0010;
	mem[1573] = 4'b0010;
	mem[1574] = 4'b0010;
	mem[1575] = 4'b0010;
	mem[1576] = 4'b0010;
	mem[1577] = 4'b0010;
	mem[1578] = 4'b0010;
	mem[1579] = 4'b0010;
	mem[1580] = 4'b0010;
	mem[1581] = 4'b0010;
	mem[1582] = 4'b0010;
	mem[1583] = 4'b0010;
	mem[1584] = 4'b0010;
	mem[1585] = 4'b0010;
	mem[1586] = 4'b0010;
	mem[1587] = 4'b0010;
	mem[1588] = 4'b0011;
	mem[1589] = 4'b0011;
	mem[1590] = 4'b0011;
	mem[1591] = 4'b0010;
	mem[1592] = 4'b0010;
	mem[1593] = 4'b0010;
	mem[1594] = 4'b0010;
	mem[1595] = 4'b0010;
	mem[1596] = 4'b0010;
	mem[1597] = 4'b0010;
	mem[1598] = 4'b0010;
	mem[1599] = 4'b0010;
	mem[1600] = 4'b0011;
	mem[1601] = 4'b0010;
	mem[1602] = 4'b0010;
	mem[1603] = 4'b0010;
	mem[1604] = 4'b0010;
	mem[1605] = 4'b0010;
	mem[1606] = 4'b0010;
	mem[1607] = 4'b1011;
	mem[1608] = 4'b1101;
	mem[1609] = 4'b1101;
	mem[1610] = 4'b1101;
	mem[1611] = 4'b1101;
	mem[1612] = 4'b1101;
	mem[1613] = 4'b1101;
	mem[1614] = 4'b1101;
	mem[1615] = 4'b1101;
	mem[1616] = 4'b1101;
	mem[1617] = 4'b1101;
	mem[1618] = 4'b1101;
	mem[1619] = 4'b1101;
	mem[1620] = 4'b1101;
	mem[1621] = 4'b1101;
	mem[1622] = 4'b1101;
	mem[1623] = 4'b1101;
	mem[1624] = 4'b0011;
	mem[1625] = 4'b0000;
	mem[1626] = 4'b0000;
	mem[1627] = 4'b0000;
	mem[1628] = 4'b0000;
	mem[1629] = 4'b0000;
	mem[1630] = 4'b0000;
	mem[1631] = 4'b0000;
	mem[1632] = 4'b0000;
	mem[1633] = 4'b0000;
	mem[1634] = 4'b0000;
	mem[1635] = 4'b0001;
	mem[1636] = 4'b0000;
	mem[1637] = 4'b0000;
	mem[1638] = 4'b0001;
	mem[1639] = 4'b0001;
	mem[1640] = 4'b0000;
	mem[1641] = 4'b0110;
	mem[1642] = 4'b1010;
	mem[1643] = 4'b1010;
	mem[1644] = 4'b1011;
	mem[1645] = 4'b1011;
	mem[1646] = 4'b1011;
	mem[1647] = 4'b1011;
	mem[1648] = 4'b1011;
	mem[1649] = 4'b1011;
	mem[1650] = 4'b1011;
	mem[1651] = 4'b1011;
	mem[1652] = 4'b1011;
	mem[1653] = 4'b1011;
	mem[1654] = 4'b1011;
	mem[1655] = 4'b1011;
	mem[1656] = 4'b1011;
	mem[1657] = 4'b1010;
	mem[1658] = 4'b0010;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0000;
	mem[1668] = 4'b0000;
	mem[1669] = 4'b0100;
	mem[1670] = 4'b0111;
	mem[1671] = 4'b0011;
	mem[1672] = 4'b0000;
	mem[1673] = 4'b0000;
	mem[1674] = 4'b0000;
	mem[1675] = 4'b0000;
	mem[1676] = 4'b0000;
	mem[1677] = 4'b0000;
	mem[1678] = 4'b0000;
	mem[1679] = 4'b0000;
	mem[1680] = 4'b0000;
	mem[1681] = 4'b0000;
	mem[1682] = 4'b0000;
	mem[1683] = 4'b0000;
	mem[1684] = 4'b0000;
	mem[1685] = 4'b0000;
	mem[1686] = 4'b0000;
	mem[1687] = 4'b0000;
	mem[1688] = 4'b0000;
	mem[1689] = 4'b0000;
	mem[1690] = 4'b0000;
	mem[1691] = 4'b0000;
	mem[1692] = 4'b0000;
	mem[1693] = 4'b0000;
	mem[1694] = 4'b0000;
	mem[1695] = 4'b0000;
	mem[1696] = 4'b0000;
	mem[1697] = 4'b0000;
	mem[1698] = 4'b0000;
	mem[1699] = 4'b0000;
	mem[1700] = 4'b0000;
	mem[1701] = 4'b0000;
	mem[1702] = 4'b0000;
	mem[1703] = 4'b0000;
	mem[1704] = 4'b0000;
	mem[1705] = 4'b0000;
	mem[1706] = 4'b0000;
	mem[1707] = 4'b0000;
	mem[1708] = 4'b0000;
	mem[1709] = 4'b0000;
	mem[1710] = 4'b0000;
	mem[1711] = 4'b0000;
	mem[1712] = 4'b0000;
	mem[1713] = 4'b0000;
	mem[1714] = 4'b0000;
	mem[1715] = 4'b0000;
	mem[1716] = 4'b0000;
	mem[1717] = 4'b0000;
	mem[1718] = 4'b0000;
	mem[1719] = 4'b0000;
	mem[1720] = 4'b0000;
	mem[1721] = 4'b0000;
	mem[1722] = 4'b0000;
	mem[1723] = 4'b0000;
	mem[1724] = 4'b0000;
	mem[1725] = 4'b0000;
	mem[1726] = 4'b0000;
	mem[1727] = 4'b0001;
	mem[1728] = 4'b0001;
	mem[1729] = 4'b0000;
	mem[1730] = 4'b0000;
	mem[1731] = 4'b0000;
	mem[1732] = 4'b0000;
	mem[1733] = 4'b0000;
	mem[1734] = 4'b0000;
	mem[1735] = 4'b1100;
	mem[1736] = 4'b1111;
	mem[1737] = 4'b1111;
	mem[1738] = 4'b1111;
	mem[1739] = 4'b1111;
	mem[1740] = 4'b1111;
	mem[1741] = 4'b1111;
	mem[1742] = 4'b1111;
	mem[1743] = 4'b1111;
	mem[1744] = 4'b1111;
	mem[1745] = 4'b1111;
	mem[1746] = 4'b1111;
	mem[1747] = 4'b1111;
	mem[1748] = 4'b1111;
	mem[1749] = 4'b1111;
	mem[1750] = 4'b1111;
	mem[1751] = 4'b1111;
	mem[1752] = 4'b0100;
	mem[1753] = 4'b0000;
	mem[1754] = 4'b0000;
	mem[1755] = 4'b0000;
	mem[1756] = 4'b0000;
	mem[1757] = 4'b0000;
	mem[1758] = 4'b0000;
	mem[1759] = 4'b0000;
	mem[1760] = 4'b0000;
	mem[1761] = 4'b0000;
	mem[1762] = 4'b0000;
	mem[1763] = 4'b0000;
	mem[1764] = 4'b0000;
	mem[1765] = 4'b0000;
	mem[1766] = 4'b0000;
	mem[1767] = 4'b0000;
	mem[1768] = 4'b0000;
	mem[1769] = 4'b0111;
	mem[1770] = 4'b1100;
	mem[1771] = 4'b1100;
	mem[1772] = 4'b1100;
	mem[1773] = 4'b1100;
	mem[1774] = 4'b1100;
	mem[1775] = 4'b1100;
	mem[1776] = 4'b1100;
	mem[1777] = 4'b1100;
	mem[1778] = 4'b1100;
	mem[1779] = 4'b1100;
	mem[1780] = 4'b1100;
	mem[1781] = 4'b1100;
	mem[1782] = 4'b1100;
	mem[1783] = 4'b1100;
	mem[1784] = 4'b1100;
	mem[1785] = 4'b1100;
	mem[1786] = 4'b0010;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0000;
	mem[1796] = 4'b0000;
	mem[1797] = 4'b0100;
	mem[1798] = 4'b0011;
	mem[1799] = 4'b0000;
	mem[1800] = 4'b0000;
	mem[1801] = 4'b0000;
	mem[1802] = 4'b0000;
	mem[1803] = 4'b0000;
	mem[1804] = 4'b0000;
	mem[1805] = 4'b0000;
	mem[1806] = 4'b0000;
	mem[1807] = 4'b0000;
	mem[1808] = 4'b0000;
	mem[1809] = 4'b0000;
	mem[1810] = 4'b0000;
	mem[1811] = 4'b0000;
	mem[1812] = 4'b0000;
	mem[1813] = 4'b0000;
	mem[1814] = 4'b0000;
	mem[1815] = 4'b0000;
	mem[1816] = 4'b0000;
	mem[1817] = 4'b0000;
	mem[1818] = 4'b0000;
	mem[1819] = 4'b0000;
	mem[1820] = 4'b0000;
	mem[1821] = 4'b0000;
	mem[1822] = 4'b0000;
	mem[1823] = 4'b0000;
	mem[1824] = 4'b0000;
	mem[1825] = 4'b0000;
	mem[1826] = 4'b0000;
	mem[1827] = 4'b0000;
	mem[1828] = 4'b0000;
	mem[1829] = 4'b0000;
	mem[1830] = 4'b0000;
	mem[1831] = 4'b0000;
	mem[1832] = 4'b0000;
	mem[1833] = 4'b0000;
	mem[1834] = 4'b0000;
	mem[1835] = 4'b0000;
	mem[1836] = 4'b0000;
	mem[1837] = 4'b0000;
	mem[1838] = 4'b0000;
	mem[1839] = 4'b0000;
	mem[1840] = 4'b0000;
	mem[1841] = 4'b0000;
	mem[1842] = 4'b0000;
	mem[1843] = 4'b0000;
	mem[1844] = 4'b0000;
	mem[1845] = 4'b0000;
	mem[1846] = 4'b0000;
	mem[1847] = 4'b0000;
	mem[1848] = 4'b0000;
	mem[1849] = 4'b0000;
	mem[1850] = 4'b0000;
	mem[1851] = 4'b0000;
	mem[1852] = 4'b0000;
	mem[1853] = 4'b0000;
	mem[1854] = 4'b0001;
	mem[1855] = 4'b0001;
	mem[1856] = 4'b0000;
	mem[1857] = 4'b0000;
	mem[1858] = 4'b0000;
	mem[1859] = 4'b0000;
	mem[1860] = 4'b0000;
	mem[1861] = 4'b0000;
	mem[1862] = 4'b0000;
	mem[1863] = 4'b1100;
	mem[1864] = 4'b1111;
	mem[1865] = 4'b1111;
	mem[1866] = 4'b1111;
	mem[1867] = 4'b1111;
	mem[1868] = 4'b1111;
	mem[1869] = 4'b1111;
	mem[1870] = 4'b1111;
	mem[1871] = 4'b1111;
	mem[1872] = 4'b1111;
	mem[1873] = 4'b1111;
	mem[1874] = 4'b1111;
	mem[1875] = 4'b1111;
	mem[1876] = 4'b1111;
	mem[1877] = 4'b1111;
	mem[1878] = 4'b1111;
	mem[1879] = 4'b1111;
	mem[1880] = 4'b0011;
	mem[1881] = 4'b0000;
	mem[1882] = 4'b0000;
	mem[1883] = 4'b0000;
	mem[1884] = 4'b0000;
	mem[1885] = 4'b0000;
	mem[1886] = 4'b0000;
	mem[1887] = 4'b0000;
	mem[1888] = 4'b0000;
	mem[1889] = 4'b0000;
	mem[1890] = 4'b0000;
	mem[1891] = 4'b0000;
	mem[1892] = 4'b0000;
	mem[1893] = 4'b0000;
	mem[1894] = 4'b0000;
	mem[1895] = 4'b0000;
	mem[1896] = 4'b0000;
	mem[1897] = 4'b0111;
	mem[1898] = 4'b1101;
	mem[1899] = 4'b1100;
	mem[1900] = 4'b1100;
	mem[1901] = 4'b1100;
	mem[1902] = 4'b1100;
	mem[1903] = 4'b1100;
	mem[1904] = 4'b1100;
	mem[1905] = 4'b1100;
	mem[1906] = 4'b1100;
	mem[1907] = 4'b1100;
	mem[1908] = 4'b1100;
	mem[1909] = 4'b1100;
	mem[1910] = 4'b1100;
	mem[1911] = 4'b1100;
	mem[1912] = 4'b1100;
	mem[1913] = 4'b1100;
	mem[1914] = 4'b0010;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0000;
	mem[1924] = 4'b0000;
	mem[1925] = 4'b0000;
	mem[1926] = 4'b0000;
	mem[1927] = 4'b0000;
	mem[1928] = 4'b0000;
	mem[1929] = 4'b0000;
	mem[1930] = 4'b0000;
	mem[1931] = 4'b0000;
	mem[1932] = 4'b0000;
	mem[1933] = 4'b0000;
	mem[1934] = 4'b0000;
	mem[1935] = 4'b0000;
	mem[1936] = 4'b0000;
	mem[1937] = 4'b0000;
	mem[1938] = 4'b0000;
	mem[1939] = 4'b0000;
	mem[1940] = 4'b0000;
	mem[1941] = 4'b0000;
	mem[1942] = 4'b0000;
	mem[1943] = 4'b0000;
	mem[1944] = 4'b0000;
	mem[1945] = 4'b0000;
	mem[1946] = 4'b0000;
	mem[1947] = 4'b0000;
	mem[1948] = 4'b0000;
	mem[1949] = 4'b0000;
	mem[1950] = 4'b0000;
	mem[1951] = 4'b0000;
	mem[1952] = 4'b0000;
	mem[1953] = 4'b0000;
	mem[1954] = 4'b0000;
	mem[1955] = 4'b0000;
	mem[1956] = 4'b0000;
	mem[1957] = 4'b0000;
	mem[1958] = 4'b0000;
	mem[1959] = 4'b0000;
	mem[1960] = 4'b0000;
	mem[1961] = 4'b0000;
	mem[1962] = 4'b0000;
	mem[1963] = 4'b0000;
	mem[1964] = 4'b0000;
	mem[1965] = 4'b0000;
	mem[1966] = 4'b0000;
	mem[1967] = 4'b0000;
	mem[1968] = 4'b0000;
	mem[1969] = 4'b0000;
	mem[1970] = 4'b0000;
	mem[1971] = 4'b0000;
	mem[1972] = 4'b0000;
	mem[1973] = 4'b0000;
	mem[1974] = 4'b0000;
	mem[1975] = 4'b0000;
	mem[1976] = 4'b0000;
	mem[1977] = 4'b0000;
	mem[1978] = 4'b0000;
	mem[1979] = 4'b0000;
	mem[1980] = 4'b0000;
	mem[1981] = 4'b0001;
	mem[1982] = 4'b0001;
	mem[1983] = 4'b0000;
	mem[1984] = 4'b0000;
	mem[1985] = 4'b0000;
	mem[1986] = 4'b0000;
	mem[1987] = 4'b0000;
	mem[1988] = 4'b0000;
	mem[1989] = 4'b0000;
	mem[1990] = 4'b0000;
	mem[1991] = 4'b1100;
	mem[1992] = 4'b1111;
	mem[1993] = 4'b1111;
	mem[1994] = 4'b1111;
	mem[1995] = 4'b1111;
	mem[1996] = 4'b1111;
	mem[1997] = 4'b1111;
	mem[1998] = 4'b1111;
	mem[1999] = 4'b1111;
	mem[2000] = 4'b1111;
	mem[2001] = 4'b1111;
	mem[2002] = 4'b1111;
	mem[2003] = 4'b1111;
	mem[2004] = 4'b1111;
	mem[2005] = 4'b1111;
	mem[2006] = 4'b1111;
	mem[2007] = 4'b1111;
	mem[2008] = 4'b0100;
	mem[2009] = 4'b0000;
	mem[2010] = 4'b0000;
	mem[2011] = 4'b0000;
	mem[2012] = 4'b0000;
	mem[2013] = 4'b0000;
	mem[2014] = 4'b0000;
	mem[2015] = 4'b0000;
	mem[2016] = 4'b0000;
	mem[2017] = 4'b0000;
	mem[2018] = 4'b0000;
	mem[2019] = 4'b0000;
	mem[2020] = 4'b0000;
	mem[2021] = 4'b0000;
	mem[2022] = 4'b0000;
	mem[2023] = 4'b0000;
	mem[2024] = 4'b0001;
	mem[2025] = 4'b1000;
	mem[2026] = 4'b1100;
	mem[2027] = 4'b1100;
	mem[2028] = 4'b1100;
	mem[2029] = 4'b1100;
	mem[2030] = 4'b1100;
	mem[2031] = 4'b1100;
	mem[2032] = 4'b1100;
	mem[2033] = 4'b1100;
	mem[2034] = 4'b1100;
	mem[2035] = 4'b1100;
	mem[2036] = 4'b1100;
	mem[2037] = 4'b1100;
	mem[2038] = 4'b1100;
	mem[2039] = 4'b1100;
	mem[2040] = 4'b1100;
	mem[2041] = 4'b1100;
	mem[2042] = 4'b0010;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0000;
	mem[2052] = 4'b0000;
	mem[2053] = 4'b0000;
	mem[2054] = 4'b0000;
	mem[2055] = 4'b0000;
	mem[2056] = 4'b0000;
	mem[2057] = 4'b0000;
	mem[2058] = 4'b0000;
	mem[2059] = 4'b0000;
	mem[2060] = 4'b0000;
	mem[2061] = 4'b0000;
	mem[2062] = 4'b0000;
	mem[2063] = 4'b0000;
	mem[2064] = 4'b0000;
	mem[2065] = 4'b0000;
	mem[2066] = 4'b0000;
	mem[2067] = 4'b0000;
	mem[2068] = 4'b0000;
	mem[2069] = 4'b0000;
	mem[2070] = 4'b0000;
	mem[2071] = 4'b0000;
	mem[2072] = 4'b0000;
	mem[2073] = 4'b0000;
	mem[2074] = 4'b0000;
	mem[2075] = 4'b0000;
	mem[2076] = 4'b0000;
	mem[2077] = 4'b0000;
	mem[2078] = 4'b0000;
	mem[2079] = 4'b0000;
	mem[2080] = 4'b0000;
	mem[2081] = 4'b0000;
	mem[2082] = 4'b0000;
	mem[2083] = 4'b0000;
	mem[2084] = 4'b0000;
	mem[2085] = 4'b0000;
	mem[2086] = 4'b0000;
	mem[2087] = 4'b0000;
	mem[2088] = 4'b0000;
	mem[2089] = 4'b0000;
	mem[2090] = 4'b0001;
	mem[2091] = 4'b0001;
	mem[2092] = 4'b0001;
	mem[2093] = 4'b0001;
	mem[2094] = 4'b0000;
	mem[2095] = 4'b0000;
	mem[2096] = 4'b0000;
	mem[2097] = 4'b0000;
	mem[2098] = 4'b0000;
	mem[2099] = 4'b0000;
	mem[2100] = 4'b0000;
	mem[2101] = 4'b0000;
	mem[2102] = 4'b0000;
	mem[2103] = 4'b0001;
	mem[2104] = 4'b0001;
	mem[2105] = 4'b0000;
	mem[2106] = 4'b0001;
	mem[2107] = 4'b0001;
	mem[2108] = 4'b0001;
	mem[2109] = 4'b0000;
	mem[2110] = 4'b0000;
	mem[2111] = 4'b0000;
	mem[2112] = 4'b0000;
	mem[2113] = 4'b0000;
	mem[2114] = 4'b0000;
	mem[2115] = 4'b0000;
	mem[2116] = 4'b0000;
	mem[2117] = 4'b0000;
	mem[2118] = 4'b0000;
	mem[2119] = 4'b1100;
	mem[2120] = 4'b1111;
	mem[2121] = 4'b1111;
	mem[2122] = 4'b1111;
	mem[2123] = 4'b1111;
	mem[2124] = 4'b1111;
	mem[2125] = 4'b1111;
	mem[2126] = 4'b1111;
	mem[2127] = 4'b1111;
	mem[2128] = 4'b1111;
	mem[2129] = 4'b1111;
	mem[2130] = 4'b1111;
	mem[2131] = 4'b1111;
	mem[2132] = 4'b1111;
	mem[2133] = 4'b1111;
	mem[2134] = 4'b1111;
	mem[2135] = 4'b1111;
	mem[2136] = 4'b0100;
	mem[2137] = 4'b0000;
	mem[2138] = 4'b0000;
	mem[2139] = 4'b0000;
	mem[2140] = 4'b0000;
	mem[2141] = 4'b0000;
	mem[2142] = 4'b0000;
	mem[2143] = 4'b0000;
	mem[2144] = 4'b0000;
	mem[2145] = 4'b0000;
	mem[2146] = 4'b0000;
	mem[2147] = 4'b0000;
	mem[2148] = 4'b0000;
	mem[2149] = 4'b0000;
	mem[2150] = 4'b0000;
	mem[2151] = 4'b0001;
	mem[2152] = 4'b0001;
	mem[2153] = 4'b1000;
	mem[2154] = 4'b1100;
	mem[2155] = 4'b1100;
	mem[2156] = 4'b1100;
	mem[2157] = 4'b1100;
	mem[2158] = 4'b1100;
	mem[2159] = 4'b1100;
	mem[2160] = 4'b1100;
	mem[2161] = 4'b1100;
	mem[2162] = 4'b1100;
	mem[2163] = 4'b1100;
	mem[2164] = 4'b1100;
	mem[2165] = 4'b1100;
	mem[2166] = 4'b1100;
	mem[2167] = 4'b1100;
	mem[2168] = 4'b1100;
	mem[2169] = 4'b1100;
	mem[2170] = 4'b0010;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0000;
	mem[2180] = 4'b0000;
	mem[2181] = 4'b0000;
	mem[2182] = 4'b0000;
	mem[2183] = 4'b0000;
	mem[2184] = 4'b0000;
	mem[2185] = 4'b0000;
	mem[2186] = 4'b0000;
	mem[2187] = 4'b0000;
	mem[2188] = 4'b0000;
	mem[2189] = 4'b0000;
	mem[2190] = 4'b0000;
	mem[2191] = 4'b0000;
	mem[2192] = 4'b0000;
	mem[2193] = 4'b0000;
	mem[2194] = 4'b0000;
	mem[2195] = 4'b0000;
	mem[2196] = 4'b0000;
	mem[2197] = 4'b0000;
	mem[2198] = 4'b0000;
	mem[2199] = 4'b0000;
	mem[2200] = 4'b0000;
	mem[2201] = 4'b0000;
	mem[2202] = 4'b0000;
	mem[2203] = 4'b0000;
	mem[2204] = 4'b0000;
	mem[2205] = 4'b0000;
	mem[2206] = 4'b0000;
	mem[2207] = 4'b0000;
	mem[2208] = 4'b0000;
	mem[2209] = 4'b0000;
	mem[2210] = 4'b0000;
	mem[2211] = 4'b0000;
	mem[2212] = 4'b0000;
	mem[2213] = 4'b0000;
	mem[2214] = 4'b0000;
	mem[2215] = 4'b0000;
	mem[2216] = 4'b0000;
	mem[2217] = 4'b0001;
	mem[2218] = 4'b0001;
	mem[2219] = 4'b0000;
	mem[2220] = 4'b0000;
	mem[2221] = 4'b0000;
	mem[2222] = 4'b0000;
	mem[2223] = 4'b0000;
	mem[2224] = 4'b0000;
	mem[2225] = 4'b0000;
	mem[2226] = 4'b0000;
	mem[2227] = 4'b0000;
	mem[2228] = 4'b0000;
	mem[2229] = 4'b0000;
	mem[2230] = 4'b0000;
	mem[2231] = 4'b0000;
	mem[2232] = 4'b0000;
	mem[2233] = 4'b0000;
	mem[2234] = 4'b0000;
	mem[2235] = 4'b0000;
	mem[2236] = 4'b0000;
	mem[2237] = 4'b0000;
	mem[2238] = 4'b0000;
	mem[2239] = 4'b0000;
	mem[2240] = 4'b0000;
	mem[2241] = 4'b0000;
	mem[2242] = 4'b0000;
	mem[2243] = 4'b0000;
	mem[2244] = 4'b0000;
	mem[2245] = 4'b0000;
	mem[2246] = 4'b0000;
	mem[2247] = 4'b1100;
	mem[2248] = 4'b1111;
	mem[2249] = 4'b1111;
	mem[2250] = 4'b1111;
	mem[2251] = 4'b1111;
	mem[2252] = 4'b1111;
	mem[2253] = 4'b1111;
	mem[2254] = 4'b1111;
	mem[2255] = 4'b1111;
	mem[2256] = 4'b1111;
	mem[2257] = 4'b1111;
	mem[2258] = 4'b1111;
	mem[2259] = 4'b1111;
	mem[2260] = 4'b1111;
	mem[2261] = 4'b1111;
	mem[2262] = 4'b1111;
	mem[2263] = 4'b1111;
	mem[2264] = 4'b0100;
	mem[2265] = 4'b0000;
	mem[2266] = 4'b0000;
	mem[2267] = 4'b0000;
	mem[2268] = 4'b0000;
	mem[2269] = 4'b0000;
	mem[2270] = 4'b0000;
	mem[2271] = 4'b0000;
	mem[2272] = 4'b0000;
	mem[2273] = 4'b0000;
	mem[2274] = 4'b0000;
	mem[2275] = 4'b0000;
	mem[2276] = 4'b0000;
	mem[2277] = 4'b0000;
	mem[2278] = 4'b0000;
	mem[2279] = 4'b0000;
	mem[2280] = 4'b0000;
	mem[2281] = 4'b1000;
	mem[2282] = 4'b1100;
	mem[2283] = 4'b1100;
	mem[2284] = 4'b1100;
	mem[2285] = 4'b1100;
	mem[2286] = 4'b1100;
	mem[2287] = 4'b1100;
	mem[2288] = 4'b1100;
	mem[2289] = 4'b1100;
	mem[2290] = 4'b1100;
	mem[2291] = 4'b1100;
	mem[2292] = 4'b1100;
	mem[2293] = 4'b1100;
	mem[2294] = 4'b1100;
	mem[2295] = 4'b1100;
	mem[2296] = 4'b1100;
	mem[2297] = 4'b1100;
	mem[2298] = 4'b0010;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0000;
	mem[2308] = 4'b0000;
	mem[2309] = 4'b0000;
	mem[2310] = 4'b0000;
	mem[2311] = 4'b0000;
	mem[2312] = 4'b0000;
	mem[2313] = 4'b0000;
	mem[2314] = 4'b0000;
	mem[2315] = 4'b0000;
	mem[2316] = 4'b0000;
	mem[2317] = 4'b0000;
	mem[2318] = 4'b0000;
	mem[2319] = 4'b0000;
	mem[2320] = 4'b0000;
	mem[2321] = 4'b0000;
	mem[2322] = 4'b0000;
	mem[2323] = 4'b0000;
	mem[2324] = 4'b0000;
	mem[2325] = 4'b0000;
	mem[2326] = 4'b0000;
	mem[2327] = 4'b0000;
	mem[2328] = 4'b0000;
	mem[2329] = 4'b0000;
	mem[2330] = 4'b0000;
	mem[2331] = 4'b0000;
	mem[2332] = 4'b0000;
	mem[2333] = 4'b0000;
	mem[2334] = 4'b0000;
	mem[2335] = 4'b0000;
	mem[2336] = 4'b0000;
	mem[2337] = 4'b0000;
	mem[2338] = 4'b0000;
	mem[2339] = 4'b0000;
	mem[2340] = 4'b0000;
	mem[2341] = 4'b0000;
	mem[2342] = 4'b0000;
	mem[2343] = 4'b0000;
	mem[2344] = 4'b0000;
	mem[2345] = 4'b0001;
	mem[2346] = 4'b0000;
	mem[2347] = 4'b0000;
	mem[2348] = 4'b0000;
	mem[2349] = 4'b0000;
	mem[2350] = 4'b0000;
	mem[2351] = 4'b0000;
	mem[2352] = 4'b0000;
	mem[2353] = 4'b0000;
	mem[2354] = 4'b0000;
	mem[2355] = 4'b0000;
	mem[2356] = 4'b0000;
	mem[2357] = 4'b0000;
	mem[2358] = 4'b0000;
	mem[2359] = 4'b0000;
	mem[2360] = 4'b0000;
	mem[2361] = 4'b0000;
	mem[2362] = 4'b0000;
	mem[2363] = 4'b0000;
	mem[2364] = 4'b0000;
	mem[2365] = 4'b0000;
	mem[2366] = 4'b0000;
	mem[2367] = 4'b0000;
	mem[2368] = 4'b0000;
	mem[2369] = 4'b0000;
	mem[2370] = 4'b0000;
	mem[2371] = 4'b0000;
	mem[2372] = 4'b0000;
	mem[2373] = 4'b0000;
	mem[2374] = 4'b0000;
	mem[2375] = 4'b1100;
	mem[2376] = 4'b1111;
	mem[2377] = 4'b1111;
	mem[2378] = 4'b1111;
	mem[2379] = 4'b1111;
	mem[2380] = 4'b1111;
	mem[2381] = 4'b1111;
	mem[2382] = 4'b1111;
	mem[2383] = 4'b1111;
	mem[2384] = 4'b1111;
	mem[2385] = 4'b1111;
	mem[2386] = 4'b1111;
	mem[2387] = 4'b1111;
	mem[2388] = 4'b1111;
	mem[2389] = 4'b1111;
	mem[2390] = 4'b1111;
	mem[2391] = 4'b1111;
	mem[2392] = 4'b0100;
	mem[2393] = 4'b0000;
	mem[2394] = 4'b0000;
	mem[2395] = 4'b0000;
	mem[2396] = 4'b0000;
	mem[2397] = 4'b0000;
	mem[2398] = 4'b0000;
	mem[2399] = 4'b0000;
	mem[2400] = 4'b0000;
	mem[2401] = 4'b0000;
	mem[2402] = 4'b0000;
	mem[2403] = 4'b0000;
	mem[2404] = 4'b0000;
	mem[2405] = 4'b0001;
	mem[2406] = 4'b0001;
	mem[2407] = 4'b0000;
	mem[2408] = 4'b0000;
	mem[2409] = 4'b1000;
	mem[2410] = 4'b1100;
	mem[2411] = 4'b1100;
	mem[2412] = 4'b1100;
	mem[2413] = 4'b1100;
	mem[2414] = 4'b1100;
	mem[2415] = 4'b1100;
	mem[2416] = 4'b1100;
	mem[2417] = 4'b1100;
	mem[2418] = 4'b1100;
	mem[2419] = 4'b1100;
	mem[2420] = 4'b1100;
	mem[2421] = 4'b1100;
	mem[2422] = 4'b1100;
	mem[2423] = 4'b1100;
	mem[2424] = 4'b1100;
	mem[2425] = 4'b1100;
	mem[2426] = 4'b0010;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0000;
	mem[2436] = 4'b0000;
	mem[2437] = 4'b0000;
	mem[2438] = 4'b0000;
	mem[2439] = 4'b0000;
	mem[2440] = 4'b0000;
	mem[2441] = 4'b0000;
	mem[2442] = 4'b0000;
	mem[2443] = 4'b0000;
	mem[2444] = 4'b0000;
	mem[2445] = 4'b0000;
	mem[2446] = 4'b0000;
	mem[2447] = 4'b0000;
	mem[2448] = 4'b0000;
	mem[2449] = 4'b0000;
	mem[2450] = 4'b0000;
	mem[2451] = 4'b0000;
	mem[2452] = 4'b0000;
	mem[2453] = 4'b0000;
	mem[2454] = 4'b0000;
	mem[2455] = 4'b0000;
	mem[2456] = 4'b0000;
	mem[2457] = 4'b0000;
	mem[2458] = 4'b0000;
	mem[2459] = 4'b0000;
	mem[2460] = 4'b0000;
	mem[2461] = 4'b0000;
	mem[2462] = 4'b0000;
	mem[2463] = 4'b0000;
	mem[2464] = 4'b0000;
	mem[2465] = 4'b0000;
	mem[2466] = 4'b0000;
	mem[2467] = 4'b0000;
	mem[2468] = 4'b0000;
	mem[2469] = 4'b0000;
	mem[2470] = 4'b0000;
	mem[2471] = 4'b0000;
	mem[2472] = 4'b0000;
	mem[2473] = 4'b0001;
	mem[2474] = 4'b0000;
	mem[2475] = 4'b0000;
	mem[2476] = 4'b0000;
	mem[2477] = 4'b0000;
	mem[2478] = 4'b0000;
	mem[2479] = 4'b0000;
	mem[2480] = 4'b0000;
	mem[2481] = 4'b0000;
	mem[2482] = 4'b0000;
	mem[2483] = 4'b0000;
	mem[2484] = 4'b0000;
	mem[2485] = 4'b0000;
	mem[2486] = 4'b0000;
	mem[2487] = 4'b0000;
	mem[2488] = 4'b0000;
	mem[2489] = 4'b0000;
	mem[2490] = 4'b0000;
	mem[2491] = 4'b0000;
	mem[2492] = 4'b0000;
	mem[2493] = 4'b0000;
	mem[2494] = 4'b0000;
	mem[2495] = 4'b0000;
	mem[2496] = 4'b0000;
	mem[2497] = 4'b0000;
	mem[2498] = 4'b0000;
	mem[2499] = 4'b0000;
	mem[2500] = 4'b0000;
	mem[2501] = 4'b0000;
	mem[2502] = 4'b0000;
	mem[2503] = 4'b1100;
	mem[2504] = 4'b1111;
	mem[2505] = 4'b1111;
	mem[2506] = 4'b1111;
	mem[2507] = 4'b1111;
	mem[2508] = 4'b1111;
	mem[2509] = 4'b1111;
	mem[2510] = 4'b1111;
	mem[2511] = 4'b1111;
	mem[2512] = 4'b1111;
	mem[2513] = 4'b1111;
	mem[2514] = 4'b1111;
	mem[2515] = 4'b1111;
	mem[2516] = 4'b1111;
	mem[2517] = 4'b1111;
	mem[2518] = 4'b1111;
	mem[2519] = 4'b1111;
	mem[2520] = 4'b0100;
	mem[2521] = 4'b0000;
	mem[2522] = 4'b0000;
	mem[2523] = 4'b0000;
	mem[2524] = 4'b0000;
	mem[2525] = 4'b0000;
	mem[2526] = 4'b0000;
	mem[2527] = 4'b0000;
	mem[2528] = 4'b0000;
	mem[2529] = 4'b0000;
	mem[2530] = 4'b0000;
	mem[2531] = 4'b0000;
	mem[2532] = 4'b0001;
	mem[2533] = 4'b0001;
	mem[2534] = 4'b0000;
	mem[2535] = 4'b0000;
	mem[2536] = 4'b0000;
	mem[2537] = 4'b1000;
	mem[2538] = 4'b1100;
	mem[2539] = 4'b1100;
	mem[2540] = 4'b1100;
	mem[2541] = 4'b1100;
	mem[2542] = 4'b1100;
	mem[2543] = 4'b1100;
	mem[2544] = 4'b1100;
	mem[2545] = 4'b1100;
	mem[2546] = 4'b1100;
	mem[2547] = 4'b1100;
	mem[2548] = 4'b1100;
	mem[2549] = 4'b1100;
	mem[2550] = 4'b1100;
	mem[2551] = 4'b1100;
	mem[2552] = 4'b1100;
	mem[2553] = 4'b1100;
	mem[2554] = 4'b0010;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b1000;
	mem[2564] = 4'b1101;
	mem[2565] = 4'b1101;
	mem[2566] = 4'b1101;
	mem[2567] = 4'b1101;
	mem[2568] = 4'b1101;
	mem[2569] = 4'b1100;
	mem[2570] = 4'b1100;
	mem[2571] = 4'b1100;
	mem[2572] = 4'b1100;
	mem[2573] = 4'b1100;
	mem[2574] = 4'b1011;
	mem[2575] = 4'b1011;
	mem[2576] = 4'b1011;
	mem[2577] = 4'b1011;
	mem[2578] = 4'b1011;
	mem[2579] = 4'b1010;
	mem[2580] = 4'b1010;
	mem[2581] = 4'b1010;
	mem[2582] = 4'b1010;
	mem[2583] = 4'b1010;
	mem[2584] = 4'b1001;
	mem[2585] = 4'b1001;
	mem[2586] = 4'b1001;
	mem[2587] = 4'b1001;
	mem[2588] = 4'b1001;
	mem[2589] = 4'b1000;
	mem[2590] = 4'b1000;
	mem[2591] = 4'b1000;
	mem[2592] = 4'b1000;
	mem[2593] = 4'b1000;
	mem[2594] = 4'b0111;
	mem[2595] = 4'b1000;
	mem[2596] = 4'b0111;
	mem[2597] = 4'b0110;
	mem[2598] = 4'b0110;
	mem[2599] = 4'b0110;
	mem[2600] = 4'b0110;
	mem[2601] = 4'b0110;
	mem[2602] = 4'b0110;
	mem[2603] = 4'b0110;
	mem[2604] = 4'b0110;
	mem[2605] = 4'b0101;
	mem[2606] = 4'b0101;
	mem[2607] = 4'b0101;
	mem[2608] = 4'b0101;
	mem[2609] = 4'b0101;
	mem[2610] = 4'b0100;
	mem[2611] = 4'b0100;
	mem[2612] = 4'b0100;
	mem[2613] = 4'b0100;
	mem[2614] = 4'b0011;
	mem[2615] = 4'b0100;
	mem[2616] = 4'b0011;
	mem[2617] = 4'b0011;
	mem[2618] = 4'b0011;
	mem[2619] = 4'b0011;
	mem[2620] = 4'b0010;
	mem[2621] = 4'b0010;
	mem[2622] = 4'b0010;
	mem[2623] = 4'b0010;
	mem[2624] = 4'b0010;
	mem[2625] = 4'b0001;
	mem[2626] = 4'b0001;
	mem[2627] = 4'b0001;
	mem[2628] = 4'b0001;
	mem[2629] = 4'b0001;
	mem[2630] = 4'b0001;
	mem[2631] = 4'b0010;
	mem[2632] = 4'b0010;
	mem[2633] = 4'b0010;
	mem[2634] = 4'b0010;
	mem[2635] = 4'b1010;
	mem[2636] = 4'b1111;
	mem[2637] = 4'b1111;
	mem[2638] = 4'b1111;
	mem[2639] = 4'b1110;
	mem[2640] = 4'b1110;
	mem[2641] = 4'b1110;
	mem[2642] = 4'b1101;
	mem[2643] = 4'b1101;
	mem[2644] = 4'b1101;
	mem[2645] = 4'b1100;
	mem[2646] = 4'b1100;
	mem[2647] = 4'b1100;
	mem[2648] = 4'b1010;
	mem[2649] = 4'b1001;
	mem[2650] = 4'b1001;
	mem[2651] = 4'b1001;
	mem[2652] = 4'b1001;
	mem[2653] = 4'b1000;
	mem[2654] = 4'b0111;
	mem[2655] = 4'b0111;
	mem[2656] = 4'b0111;
	mem[2657] = 4'b0110;
	mem[2658] = 4'b0110;
	mem[2659] = 4'b0111;
	mem[2660] = 4'b0111;
	mem[2661] = 4'b0110;
	mem[2662] = 4'b0101;
	mem[2663] = 4'b0101;
	mem[2664] = 4'b0101;
	mem[2665] = 4'b0110;
	mem[2666] = 4'b0110;
	mem[2667] = 4'b0110;
	mem[2668] = 4'b0101;
	mem[2669] = 4'b0101;
	mem[2670] = 4'b0101;
	mem[2671] = 4'b0101;
	mem[2672] = 4'b0100;
	mem[2673] = 4'b0100;
	mem[2674] = 4'b0100;
	mem[2675] = 4'b0100;
	mem[2676] = 4'b0011;
	mem[2677] = 4'b0011;
	mem[2678] = 4'b0011;
	mem[2679] = 4'b0011;
	mem[2680] = 4'b0011;
	mem[2681] = 4'b0010;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b1001;
	mem[2692] = 4'b1111;
	mem[2693] = 4'b1111;
	mem[2694] = 4'b1111;
	mem[2695] = 4'b1111;
	mem[2696] = 4'b1110;
	mem[2697] = 4'b1110;
	mem[2698] = 4'b1110;
	mem[2699] = 4'b1110;
	mem[2700] = 4'b1101;
	mem[2701] = 4'b1101;
	mem[2702] = 4'b1101;
	mem[2703] = 4'b1101;
	mem[2704] = 4'b1101;
	mem[2705] = 4'b1100;
	mem[2706] = 4'b1100;
	mem[2707] = 4'b1100;
	mem[2708] = 4'b1100;
	mem[2709] = 4'b1011;
	mem[2710] = 4'b1011;
	mem[2711] = 4'b1011;
	mem[2712] = 4'b1011;
	mem[2713] = 4'b1011;
	mem[2714] = 4'b1010;
	mem[2715] = 4'b1010;
	mem[2716] = 4'b1010;
	mem[2717] = 4'b1010;
	mem[2718] = 4'b1001;
	mem[2719] = 4'b1001;
	mem[2720] = 4'b1001;
	mem[2721] = 4'b1001;
	mem[2722] = 4'b1001;
	mem[2723] = 4'b1000;
	mem[2724] = 4'b1000;
	mem[2725] = 4'b0111;
	mem[2726] = 4'b0111;
	mem[2727] = 4'b0111;
	mem[2728] = 4'b0111;
	mem[2729] = 4'b0110;
	mem[2730] = 4'b0111;
	mem[2731] = 4'b0111;
	mem[2732] = 4'b0110;
	mem[2733] = 4'b0110;
	mem[2734] = 4'b0110;
	mem[2735] = 4'b0110;
	mem[2736] = 4'b0101;
	mem[2737] = 4'b0101;
	mem[2738] = 4'b0101;
	mem[2739] = 4'b0100;
	mem[2740] = 4'b0100;
	mem[2741] = 4'b0100;
	mem[2742] = 4'b0100;
	mem[2743] = 4'b0101;
	mem[2744] = 4'b0100;
	mem[2745] = 4'b0100;
	mem[2746] = 4'b0011;
	mem[2747] = 4'b0011;
	mem[2748] = 4'b0011;
	mem[2749] = 4'b0011;
	mem[2750] = 4'b0010;
	mem[2751] = 4'b0010;
	mem[2752] = 4'b0010;
	mem[2753] = 4'b0010;
	mem[2754] = 4'b0010;
	mem[2755] = 4'b0001;
	mem[2756] = 4'b0001;
	mem[2757] = 4'b0001;
	mem[2758] = 4'b0001;
	mem[2759] = 4'b0000;
	mem[2760] = 4'b0000;
	mem[2761] = 4'b0000;
	mem[2762] = 4'b0000;
	mem[2763] = 4'b1001;
	mem[2764] = 4'b1111;
	mem[2765] = 4'b1111;
	mem[2766] = 4'b1110;
	mem[2767] = 4'b1110;
	mem[2768] = 4'b1110;
	mem[2769] = 4'b1101;
	mem[2770] = 4'b1101;
	mem[2771] = 4'b1101;
	mem[2772] = 4'b1100;
	mem[2773] = 4'b1100;
	mem[2774] = 4'b1100;
	mem[2775] = 4'b1011;
	mem[2776] = 4'b1011;
	mem[2777] = 4'b1011;
	mem[2778] = 4'b1010;
	mem[2779] = 4'b1001;
	mem[2780] = 4'b1010;
	mem[2781] = 4'b1001;
	mem[2782] = 4'b1001;
	mem[2783] = 4'b1000;
	mem[2784] = 4'b0111;
	mem[2785] = 4'b0111;
	mem[2786] = 4'b1000;
	mem[2787] = 4'b1000;
	mem[2788] = 4'b0111;
	mem[2789] = 4'b0111;
	mem[2790] = 4'b0110;
	mem[2791] = 4'b0110;
	mem[2792] = 4'b0110;
	mem[2793] = 4'b0101;
	mem[2794] = 4'b0101;
	mem[2795] = 4'b0101;
	mem[2796] = 4'b0100;
	mem[2797] = 4'b0100;
	mem[2798] = 4'b0100;
	mem[2799] = 4'b0100;
	mem[2800] = 4'b0011;
	mem[2801] = 4'b0011;
	mem[2802] = 4'b0011;
	mem[2803] = 4'b0011;
	mem[2804] = 4'b0010;
	mem[2805] = 4'b0010;
	mem[2806] = 4'b0010;
	mem[2807] = 4'b0010;
	mem[2808] = 4'b0010;
	mem[2809] = 4'b0001;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b1001;
	mem[2820] = 4'b1111;
	mem[2821] = 4'b1111;
	mem[2822] = 4'b1111;
	mem[2823] = 4'b1111;
	mem[2824] = 4'b1110;
	mem[2825] = 4'b1110;
	mem[2826] = 4'b1110;
	mem[2827] = 4'b1110;
	mem[2828] = 4'b1101;
	mem[2829] = 4'b1101;
	mem[2830] = 4'b1101;
	mem[2831] = 4'b1101;
	mem[2832] = 4'b1101;
	mem[2833] = 4'b1100;
	mem[2834] = 4'b1100;
	mem[2835] = 4'b1100;
	mem[2836] = 4'b1100;
	mem[2837] = 4'b1011;
	mem[2838] = 4'b1011;
	mem[2839] = 4'b1011;
	mem[2840] = 4'b1011;
	mem[2841] = 4'b1011;
	mem[2842] = 4'b1010;
	mem[2843] = 4'b1010;
	mem[2844] = 4'b1010;
	mem[2845] = 4'b1010;
	mem[2846] = 4'b1001;
	mem[2847] = 4'b1001;
	mem[2848] = 4'b1001;
	mem[2849] = 4'b1001;
	mem[2850] = 4'b1001;
	mem[2851] = 4'b1000;
	mem[2852] = 4'b1000;
	mem[2853] = 4'b1000;
	mem[2854] = 4'b0111;
	mem[2855] = 4'b0111;
	mem[2856] = 4'b0111;
	mem[2857] = 4'b0110;
	mem[2858] = 4'b0110;
	mem[2859] = 4'b0111;
	mem[2860] = 4'b0111;
	mem[2861] = 4'b0110;
	mem[2862] = 4'b0110;
	mem[2863] = 4'b0110;
	mem[2864] = 4'b0101;
	mem[2865] = 4'b0101;
	mem[2866] = 4'b0101;
	mem[2867] = 4'b0101;
	mem[2868] = 4'b0100;
	mem[2869] = 4'b0100;
	mem[2870] = 4'b0101;
	mem[2871] = 4'b0100;
	mem[2872] = 4'b0100;
	mem[2873] = 4'b0100;
	mem[2874] = 4'b0011;
	mem[2875] = 4'b0011;
	mem[2876] = 4'b0011;
	mem[2877] = 4'b0011;
	mem[2878] = 4'b0010;
	mem[2879] = 4'b0010;
	mem[2880] = 4'b0010;
	mem[2881] = 4'b0010;
	mem[2882] = 4'b0010;
	mem[2883] = 4'b0001;
	mem[2884] = 4'b0001;
	mem[2885] = 4'b0001;
	mem[2886] = 4'b0001;
	mem[2887] = 4'b0000;
	mem[2888] = 4'b0000;
	mem[2889] = 4'b0000;
	mem[2890] = 4'b0000;
	mem[2891] = 4'b1001;
	mem[2892] = 4'b1111;
	mem[2893] = 4'b1111;
	mem[2894] = 4'b1110;
	mem[2895] = 4'b1110;
	mem[2896] = 4'b1110;
	mem[2897] = 4'b1101;
	mem[2898] = 4'b1101;
	mem[2899] = 4'b1101;
	mem[2900] = 4'b1100;
	mem[2901] = 4'b1100;
	mem[2902] = 4'b1100;
	mem[2903] = 4'b1011;
	mem[2904] = 4'b1011;
	mem[2905] = 4'b1010;
	mem[2906] = 4'b1001;
	mem[2907] = 4'b1001;
	mem[2908] = 4'b1001;
	mem[2909] = 4'b1010;
	mem[2910] = 4'b1001;
	mem[2911] = 4'b1000;
	mem[2912] = 4'b0111;
	mem[2913] = 4'b1000;
	mem[2914] = 4'b1000;
	mem[2915] = 4'b0111;
	mem[2916] = 4'b0111;
	mem[2917] = 4'b0111;
	mem[2918] = 4'b0110;
	mem[2919] = 4'b0110;
	mem[2920] = 4'b0110;
	mem[2921] = 4'b0101;
	mem[2922] = 4'b0101;
	mem[2923] = 4'b0101;
	mem[2924] = 4'b0101;
	mem[2925] = 4'b0100;
	mem[2926] = 4'b0100;
	mem[2927] = 4'b0100;
	mem[2928] = 4'b0100;
	mem[2929] = 4'b0011;
	mem[2930] = 4'b0011;
	mem[2931] = 4'b0011;
	mem[2932] = 4'b0011;
	mem[2933] = 4'b0010;
	mem[2934] = 4'b0010;
	mem[2935] = 4'b0010;
	mem[2936] = 4'b0010;
	mem[2937] = 4'b0010;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b1001;
	mem[2948] = 4'b1111;
	mem[2949] = 4'b1111;
	mem[2950] = 4'b1111;
	mem[2951] = 4'b1111;
	mem[2952] = 4'b1110;
	mem[2953] = 4'b1110;
	mem[2954] = 4'b1110;
	mem[2955] = 4'b1110;
	mem[2956] = 4'b1101;
	mem[2957] = 4'b1101;
	mem[2958] = 4'b1101;
	mem[2959] = 4'b1101;
	mem[2960] = 4'b1101;
	mem[2961] = 4'b1100;
	mem[2962] = 4'b1100;
	mem[2963] = 4'b1100;
	mem[2964] = 4'b1100;
	mem[2965] = 4'b1011;
	mem[2966] = 4'b1011;
	mem[2967] = 4'b1011;
	mem[2968] = 4'b1011;
	mem[2969] = 4'b1011;
	mem[2970] = 4'b1010;
	mem[2971] = 4'b1010;
	mem[2972] = 4'b1010;
	mem[2973] = 4'b1010;
	mem[2974] = 4'b1001;
	mem[2975] = 4'b1001;
	mem[2976] = 4'b1001;
	mem[2977] = 4'b1001;
	mem[2978] = 4'b1001;
	mem[2979] = 4'b1000;
	mem[2980] = 4'b1000;
	mem[2981] = 4'b1000;
	mem[2982] = 4'b1000;
	mem[2983] = 4'b0111;
	mem[2984] = 4'b0110;
	mem[2985] = 4'b0110;
	mem[2986] = 4'b0110;
	mem[2987] = 4'b0110;
	mem[2988] = 4'b0111;
	mem[2989] = 4'b0110;
	mem[2990] = 4'b0110;
	mem[2991] = 4'b0110;
	mem[2992] = 4'b0101;
	mem[2993] = 4'b0101;
	mem[2994] = 4'b0101;
	mem[2995] = 4'b0101;
	mem[2996] = 4'b0101;
	mem[2997] = 4'b0101;
	mem[2998] = 4'b0101;
	mem[2999] = 4'b0100;
	mem[3000] = 4'b0100;
	mem[3001] = 4'b0100;
	mem[3002] = 4'b0011;
	mem[3003] = 4'b0011;
	mem[3004] = 4'b0011;
	mem[3005] = 4'b0011;
	mem[3006] = 4'b0010;
	mem[3007] = 4'b0010;
	mem[3008] = 4'b0010;
	mem[3009] = 4'b0010;
	mem[3010] = 4'b0010;
	mem[3011] = 4'b0001;
	mem[3012] = 4'b0001;
	mem[3013] = 4'b0001;
	mem[3014] = 4'b0001;
	mem[3015] = 4'b0000;
	mem[3016] = 4'b0000;
	mem[3017] = 4'b0000;
	mem[3018] = 4'b0000;
	mem[3019] = 4'b1001;
	mem[3020] = 4'b1111;
	mem[3021] = 4'b1111;
	mem[3022] = 4'b1110;
	mem[3023] = 4'b1110;
	mem[3024] = 4'b1110;
	mem[3025] = 4'b1101;
	mem[3026] = 4'b1101;
	mem[3027] = 4'b1101;
	mem[3028] = 4'b1100;
	mem[3029] = 4'b1100;
	mem[3030] = 4'b1100;
	mem[3031] = 4'b1011;
	mem[3032] = 4'b1010;
	mem[3033] = 4'b1001;
	mem[3034] = 4'b1001;
	mem[3035] = 4'b1001;
	mem[3036] = 4'b1010;
	mem[3037] = 4'b1010;
	mem[3038] = 4'b1001;
	mem[3039] = 4'b1001;
	mem[3040] = 4'b1001;
	mem[3041] = 4'b1001;
	mem[3042] = 4'b1000;
	mem[3043] = 4'b0111;
	mem[3044] = 4'b0111;
	mem[3045] = 4'b0111;
	mem[3046] = 4'b0110;
	mem[3047] = 4'b0110;
	mem[3048] = 4'b0110;
	mem[3049] = 4'b0110;
	mem[3050] = 4'b0101;
	mem[3051] = 4'b0101;
	mem[3052] = 4'b0101;
	mem[3053] = 4'b0101;
	mem[3054] = 4'b0100;
	mem[3055] = 4'b0100;
	mem[3056] = 4'b0100;
	mem[3057] = 4'b0100;
	mem[3058] = 4'b0011;
	mem[3059] = 4'b0011;
	mem[3060] = 4'b0011;
	mem[3061] = 4'b0011;
	mem[3062] = 4'b0011;
	mem[3063] = 4'b0010;
	mem[3064] = 4'b0010;
	mem[3065] = 4'b0010;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b1001;
	mem[3076] = 4'b1111;
	mem[3077] = 4'b1111;
	mem[3078] = 4'b1111;
	mem[3079] = 4'b1111;
	mem[3080] = 4'b1110;
	mem[3081] = 4'b1110;
	mem[3082] = 4'b1110;
	mem[3083] = 4'b1110;
	mem[3084] = 4'b1101;
	mem[3085] = 4'b1101;
	mem[3086] = 4'b1101;
	mem[3087] = 4'b1101;
	mem[3088] = 4'b1101;
	mem[3089] = 4'b1100;
	mem[3090] = 4'b1100;
	mem[3091] = 4'b1100;
	mem[3092] = 4'b1100;
	mem[3093] = 4'b1011;
	mem[3094] = 4'b1011;
	mem[3095] = 4'b1011;
	mem[3096] = 4'b1011;
	mem[3097] = 4'b1011;
	mem[3098] = 4'b1010;
	mem[3099] = 4'b1010;
	mem[3100] = 4'b1010;
	mem[3101] = 4'b1010;
	mem[3102] = 4'b1001;
	mem[3103] = 4'b1001;
	mem[3104] = 4'b1001;
	mem[3105] = 4'b1001;
	mem[3106] = 4'b1001;
	mem[3107] = 4'b1000;
	mem[3108] = 4'b1000;
	mem[3109] = 4'b1000;
	mem[3110] = 4'b1000;
	mem[3111] = 4'b1000;
	mem[3112] = 4'b0111;
	mem[3113] = 4'b0110;
	mem[3114] = 4'b0110;
	mem[3115] = 4'b0110;
	mem[3116] = 4'b0110;
	mem[3117] = 4'b0110;
	mem[3118] = 4'b0110;
	mem[3119] = 4'b0110;
	mem[3120] = 4'b0101;
	mem[3121] = 4'b0101;
	mem[3122] = 4'b0101;
	mem[3123] = 4'b0101;
	mem[3124] = 4'b0101;
	mem[3125] = 4'b0101;
	mem[3126] = 4'b0100;
	mem[3127] = 4'b0100;
	mem[3128] = 4'b0100;
	mem[3129] = 4'b0100;
	mem[3130] = 4'b0011;
	mem[3131] = 4'b0011;
	mem[3132] = 4'b0011;
	mem[3133] = 4'b0011;
	mem[3134] = 4'b0010;
	mem[3135] = 4'b0010;
	mem[3136] = 4'b0010;
	mem[3137] = 4'b0010;
	mem[3138] = 4'b0010;
	mem[3139] = 4'b0001;
	mem[3140] = 4'b0001;
	mem[3141] = 4'b0001;
	mem[3142] = 4'b0001;
	mem[3143] = 4'b0000;
	mem[3144] = 4'b0000;
	mem[3145] = 4'b0000;
	mem[3146] = 4'b0000;
	mem[3147] = 4'b1001;
	mem[3148] = 4'b1111;
	mem[3149] = 4'b1111;
	mem[3150] = 4'b1110;
	mem[3151] = 4'b1110;
	mem[3152] = 4'b1110;
	mem[3153] = 4'b1101;
	mem[3154] = 4'b1101;
	mem[3155] = 4'b1100;
	mem[3156] = 4'b1011;
	mem[3157] = 4'b1011;
	mem[3158] = 4'b1100;
	mem[3159] = 4'b1011;
	mem[3160] = 4'b1011;
	mem[3161] = 4'b1001;
	mem[3162] = 4'b1001;
	mem[3163] = 4'b1011;
	mem[3164] = 4'b1010;
	mem[3165] = 4'b1001;
	mem[3166] = 4'b1001;
	mem[3167] = 4'b1001;
	mem[3168] = 4'b1000;
	mem[3169] = 4'b1000;
	mem[3170] = 4'b1000;
	mem[3171] = 4'b0111;
	mem[3172] = 4'b0111;
	mem[3173] = 4'b0111;
	mem[3174] = 4'b0110;
	mem[3175] = 4'b0110;
	mem[3176] = 4'b0110;
	mem[3177] = 4'b0110;
	mem[3178] = 4'b0101;
	mem[3179] = 4'b0101;
	mem[3180] = 4'b0101;
	mem[3181] = 4'b0101;
	mem[3182] = 4'b0100;
	mem[3183] = 4'b0100;
	mem[3184] = 4'b0100;
	mem[3185] = 4'b0100;
	mem[3186] = 4'b0100;
	mem[3187] = 4'b0011;
	mem[3188] = 4'b0011;
	mem[3189] = 4'b0011;
	mem[3190] = 4'b0011;
	mem[3191] = 4'b0011;
	mem[3192] = 4'b0010;
	mem[3193] = 4'b0010;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b1001;
	mem[3204] = 4'b1111;
	mem[3205] = 4'b1111;
	mem[3206] = 4'b1111;
	mem[3207] = 4'b1111;
	mem[3208] = 4'b1110;
	mem[3209] = 4'b1110;
	mem[3210] = 4'b1110;
	mem[3211] = 4'b1110;
	mem[3212] = 4'b1101;
	mem[3213] = 4'b1101;
	mem[3214] = 4'b1101;
	mem[3215] = 4'b1101;
	mem[3216] = 4'b1101;
	mem[3217] = 4'b1100;
	mem[3218] = 4'b1100;
	mem[3219] = 4'b1100;
	mem[3220] = 4'b1100;
	mem[3221] = 4'b1011;
	mem[3222] = 4'b1011;
	mem[3223] = 4'b1011;
	mem[3224] = 4'b1011;
	mem[3225] = 4'b1011;
	mem[3226] = 4'b1010;
	mem[3227] = 4'b1010;
	mem[3228] = 4'b1010;
	mem[3229] = 4'b1001;
	mem[3230] = 4'b1001;
	mem[3231] = 4'b1000;
	mem[3232] = 4'b1000;
	mem[3233] = 4'b1000;
	mem[3234] = 4'b1000;
	mem[3235] = 4'b1000;
	mem[3236] = 4'b1000;
	mem[3237] = 4'b1000;
	mem[3238] = 4'b1000;
	mem[3239] = 4'b0111;
	mem[3240] = 4'b1000;
	mem[3241] = 4'b0110;
	mem[3242] = 4'b0110;
	mem[3243] = 4'b0110;
	mem[3244] = 4'b0110;
	mem[3245] = 4'b0101;
	mem[3246] = 4'b0110;
	mem[3247] = 4'b0110;
	mem[3248] = 4'b0101;
	mem[3249] = 4'b0101;
	mem[3250] = 4'b0101;
	mem[3251] = 4'b0101;
	mem[3252] = 4'b0101;
	mem[3253] = 4'b0100;
	mem[3254] = 4'b0100;
	mem[3255] = 4'b0100;
	mem[3256] = 4'b0100;
	mem[3257] = 4'b0100;
	mem[3258] = 4'b0011;
	mem[3259] = 4'b0011;
	mem[3260] = 4'b0011;
	mem[3261] = 4'b0011;
	mem[3262] = 4'b0010;
	mem[3263] = 4'b0010;
	mem[3264] = 4'b0010;
	mem[3265] = 4'b0010;
	mem[3266] = 4'b0010;
	mem[3267] = 4'b0001;
	mem[3268] = 4'b0001;
	mem[3269] = 4'b0001;
	mem[3270] = 4'b0001;
	mem[3271] = 4'b0000;
	mem[3272] = 4'b0000;
	mem[3273] = 4'b0000;
	mem[3274] = 4'b0000;
	mem[3275] = 4'b1001;
	mem[3276] = 4'b1111;
	mem[3277] = 4'b1111;
	mem[3278] = 4'b1110;
	mem[3279] = 4'b1110;
	mem[3280] = 4'b1110;
	mem[3281] = 4'b1101;
	mem[3282] = 4'b1100;
	mem[3283] = 4'b1011;
	mem[3284] = 4'b1011;
	mem[3285] = 4'b1100;
	mem[3286] = 4'b1100;
	mem[3287] = 4'b1011;
	mem[3288] = 4'b1011;
	mem[3289] = 4'b1011;
	mem[3290] = 4'b1011;
	mem[3291] = 4'b1010;
	mem[3292] = 4'b1010;
	mem[3293] = 4'b1001;
	mem[3294] = 4'b1001;
	mem[3295] = 4'b1001;
	mem[3296] = 4'b1000;
	mem[3297] = 4'b1000;
	mem[3298] = 4'b1000;
	mem[3299] = 4'b0111;
	mem[3300] = 4'b0111;
	mem[3301] = 4'b0111;
	mem[3302] = 4'b0111;
	mem[3303] = 4'b0110;
	mem[3304] = 4'b0110;
	mem[3305] = 4'b0110;
	mem[3306] = 4'b0110;
	mem[3307] = 4'b0101;
	mem[3308] = 4'b0101;
	mem[3309] = 4'b0101;
	mem[3310] = 4'b0101;
	mem[3311] = 4'b0100;
	mem[3312] = 4'b0100;
	mem[3313] = 4'b0100;
	mem[3314] = 4'b0100;
	mem[3315] = 4'b0100;
	mem[3316] = 4'b0011;
	mem[3317] = 4'b0011;
	mem[3318] = 4'b0011;
	mem[3319] = 4'b0011;
	mem[3320] = 4'b0011;
	mem[3321] = 4'b0010;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b1001;
	mem[3332] = 4'b1111;
	mem[3333] = 4'b1111;
	mem[3334] = 4'b1111;
	mem[3335] = 4'b1111;
	mem[3336] = 4'b1110;
	mem[3337] = 4'b1110;
	mem[3338] = 4'b1110;
	mem[3339] = 4'b1110;
	mem[3340] = 4'b1101;
	mem[3341] = 4'b1101;
	mem[3342] = 4'b1101;
	mem[3343] = 4'b1101;
	mem[3344] = 4'b1101;
	mem[3345] = 4'b1100;
	mem[3346] = 4'b1100;
	mem[3347] = 4'b1100;
	mem[3348] = 4'b1100;
	mem[3349] = 4'b1011;
	mem[3350] = 4'b1011;
	mem[3351] = 4'b1011;
	mem[3352] = 4'b1011;
	mem[3353] = 4'b1011;
	mem[3354] = 4'b1010;
	mem[3355] = 4'b1010;
	mem[3356] = 4'b1001;
	mem[3357] = 4'b1001;
	mem[3358] = 4'b1000;
	mem[3359] = 4'b1000;
	mem[3360] = 4'b1000;
	mem[3361] = 4'b1000;
	mem[3362] = 4'b1000;
	mem[3363] = 4'b0111;
	mem[3364] = 4'b0111;
	mem[3365] = 4'b1000;
	mem[3366] = 4'b1000;
	mem[3367] = 4'b0111;
	mem[3368] = 4'b0111;
	mem[3369] = 4'b0111;
	mem[3370] = 4'b0110;
	mem[3371] = 4'b0110;
	mem[3372] = 4'b0110;
	mem[3373] = 4'b0110;
	mem[3374] = 4'b0101;
	mem[3375] = 4'b0110;
	mem[3376] = 4'b0110;
	mem[3377] = 4'b0101;
	mem[3378] = 4'b0101;
	mem[3379] = 4'b0101;
	mem[3380] = 4'b0101;
	mem[3381] = 4'b0100;
	mem[3382] = 4'b0100;
	mem[3383] = 4'b0100;
	mem[3384] = 4'b0100;
	mem[3385] = 4'b0100;
	mem[3386] = 4'b0011;
	mem[3387] = 4'b0011;
	mem[3388] = 4'b0011;
	mem[3389] = 4'b0011;
	mem[3390] = 4'b0010;
	mem[3391] = 4'b0010;
	mem[3392] = 4'b0010;
	mem[3393] = 4'b0010;
	mem[3394] = 4'b0010;
	mem[3395] = 4'b0001;
	mem[3396] = 4'b0001;
	mem[3397] = 4'b0001;
	mem[3398] = 4'b0001;
	mem[3399] = 4'b0000;
	mem[3400] = 4'b0000;
	mem[3401] = 4'b0000;
	mem[3402] = 4'b0000;
	mem[3403] = 4'b1001;
	mem[3404] = 4'b1111;
	mem[3405] = 4'b1111;
	mem[3406] = 4'b1110;
	mem[3407] = 4'b1110;
	mem[3408] = 4'b1110;
	mem[3409] = 4'b1100;
	mem[3410] = 4'b1011;
	mem[3411] = 4'b1100;
	mem[3412] = 4'b1100;
	mem[3413] = 4'b1100;
	mem[3414] = 4'b1011;
	mem[3415] = 4'b1010;
	mem[3416] = 4'b1011;
	mem[3417] = 4'b1011;
	mem[3418] = 4'b1010;
	mem[3419] = 4'b1010;
	mem[3420] = 4'b1010;
	mem[3421] = 4'b1001;
	mem[3422] = 4'b1001;
	mem[3423] = 4'b1001;
	mem[3424] = 4'b1000;
	mem[3425] = 4'b1000;
	mem[3426] = 4'b1000;
	mem[3427] = 4'b1000;
	mem[3428] = 4'b0111;
	mem[3429] = 4'b0111;
	mem[3430] = 4'b0111;
	mem[3431] = 4'b0111;
	mem[3432] = 4'b0110;
	mem[3433] = 4'b0110;
	mem[3434] = 4'b0110;
	mem[3435] = 4'b0110;
	mem[3436] = 4'b0101;
	mem[3437] = 4'b0101;
	mem[3438] = 4'b0101;
	mem[3439] = 4'b0101;
	mem[3440] = 4'b0100;
	mem[3441] = 4'b0100;
	mem[3442] = 4'b0100;
	mem[3443] = 4'b0100;
	mem[3444] = 4'b0100;
	mem[3445] = 4'b0011;
	mem[3446] = 4'b0011;
	mem[3447] = 4'b0011;
	mem[3448] = 4'b0011;
	mem[3449] = 4'b0011;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b1001;
	mem[3460] = 4'b1111;
	mem[3461] = 4'b1111;
	mem[3462] = 4'b1111;
	mem[3463] = 4'b1111;
	mem[3464] = 4'b1110;
	mem[3465] = 4'b1110;
	mem[3466] = 4'b1110;
	mem[3467] = 4'b1110;
	mem[3468] = 4'b1101;
	mem[3469] = 4'b1101;
	mem[3470] = 4'b1101;
	mem[3471] = 4'b1101;
	mem[3472] = 4'b1101;
	mem[3473] = 4'b1100;
	mem[3474] = 4'b1100;
	mem[3475] = 4'b1100;
	mem[3476] = 4'b1100;
	mem[3477] = 4'b1011;
	mem[3478] = 4'b1011;
	mem[3479] = 4'b1011;
	mem[3480] = 4'b1011;
	mem[3481] = 4'b1011;
	mem[3482] = 4'b1010;
	mem[3483] = 4'b1001;
	mem[3484] = 4'b1001;
	mem[3485] = 4'b1001;
	mem[3486] = 4'b1000;
	mem[3487] = 4'b1000;
	mem[3488] = 4'b1000;
	mem[3489] = 4'b1000;
	mem[3490] = 4'b1000;
	mem[3491] = 4'b0111;
	mem[3492] = 4'b0111;
	mem[3493] = 4'b0111;
	mem[3494] = 4'b1000;
	mem[3495] = 4'b1000;
	mem[3496] = 4'b0111;
	mem[3497] = 4'b0111;
	mem[3498] = 4'b0111;
	mem[3499] = 4'b0110;
	mem[3500] = 4'b0110;
	mem[3501] = 4'b0110;
	mem[3502] = 4'b0101;
	mem[3503] = 4'b0101;
	mem[3504] = 4'b0110;
	mem[3505] = 4'b0101;
	mem[3506] = 4'b0101;
	mem[3507] = 4'b0101;
	mem[3508] = 4'b0101;
	mem[3509] = 4'b0100;
	mem[3510] = 4'b0100;
	mem[3511] = 4'b0100;
	mem[3512] = 4'b0100;
	mem[3513] = 4'b0100;
	mem[3514] = 4'b0011;
	mem[3515] = 4'b0011;
	mem[3516] = 4'b0011;
	mem[3517] = 4'b0011;
	mem[3518] = 4'b0010;
	mem[3519] = 4'b0010;
	mem[3520] = 4'b0010;
	mem[3521] = 4'b0010;
	mem[3522] = 4'b0010;
	mem[3523] = 4'b0001;
	mem[3524] = 4'b0001;
	mem[3525] = 4'b0001;
	mem[3526] = 4'b0001;
	mem[3527] = 4'b0000;
	mem[3528] = 4'b0000;
	mem[3529] = 4'b0000;
	mem[3530] = 4'b0000;
	mem[3531] = 4'b1001;
	mem[3532] = 4'b1111;
	mem[3533] = 4'b1111;
	mem[3534] = 4'b1110;
	mem[3535] = 4'b1110;
	mem[3536] = 4'b1101;
	mem[3537] = 4'b1100;
	mem[3538] = 4'b1101;
	mem[3539] = 4'b1101;
	mem[3540] = 4'b1100;
	mem[3541] = 4'b1011;
	mem[3542] = 4'b1010;
	mem[3543] = 4'b1010;
	mem[3544] = 4'b1001;
	mem[3545] = 4'b1011;
	mem[3546] = 4'b1010;
	mem[3547] = 4'b1010;
	mem[3548] = 4'b1010;
	mem[3549] = 4'b1001;
	mem[3550] = 4'b1001;
	mem[3551] = 4'b1001;
	mem[3552] = 4'b1001;
	mem[3553] = 4'b1000;
	mem[3554] = 4'b1000;
	mem[3555] = 4'b1000;
	mem[3556] = 4'b0111;
	mem[3557] = 4'b0111;
	mem[3558] = 4'b0111;
	mem[3559] = 4'b0111;
	mem[3560] = 4'b0110;
	mem[3561] = 4'b0110;
	mem[3562] = 4'b0110;
	mem[3563] = 4'b0110;
	mem[3564] = 4'b0110;
	mem[3565] = 4'b0101;
	mem[3566] = 4'b0101;
	mem[3567] = 4'b0101;
	mem[3568] = 4'b0101;
	mem[3569] = 4'b0100;
	mem[3570] = 4'b0100;
	mem[3571] = 4'b0100;
	mem[3572] = 4'b0100;
	mem[3573] = 4'b0100;
	mem[3574] = 4'b0100;
	mem[3575] = 4'b0011;
	mem[3576] = 4'b0011;
	mem[3577] = 4'b0011;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b1001;
	mem[3588] = 4'b1111;
	mem[3589] = 4'b1111;
	mem[3590] = 4'b1111;
	mem[3591] = 4'b1111;
	mem[3592] = 4'b1110;
	mem[3593] = 4'b1110;
	mem[3594] = 4'b1110;
	mem[3595] = 4'b1110;
	mem[3596] = 4'b1101;
	mem[3597] = 4'b1101;
	mem[3598] = 4'b1101;
	mem[3599] = 4'b1101;
	mem[3600] = 4'b1101;
	mem[3601] = 4'b1100;
	mem[3602] = 4'b1100;
	mem[3603] = 4'b1100;
	mem[3604] = 4'b1100;
	mem[3605] = 4'b1011;
	mem[3606] = 4'b1011;
	mem[3607] = 4'b1011;
	mem[3608] = 4'b1011;
	mem[3609] = 4'b1011;
	mem[3610] = 4'b1010;
	mem[3611] = 4'b1001;
	mem[3612] = 4'b1001;
	mem[3613] = 4'b1001;
	mem[3614] = 4'b1001;
	mem[3615] = 4'b1001;
	mem[3616] = 4'b1001;
	mem[3617] = 4'b1000;
	mem[3618] = 4'b1000;
	mem[3619] = 4'b0111;
	mem[3620] = 4'b0111;
	mem[3621] = 4'b0111;
	mem[3622] = 4'b0111;
	mem[3623] = 4'b1000;
	mem[3624] = 4'b0111;
	mem[3625] = 4'b0111;
	mem[3626] = 4'b0111;
	mem[3627] = 4'b0111;
	mem[3628] = 4'b0110;
	mem[3629] = 4'b0110;
	mem[3630] = 4'b0101;
	mem[3631] = 4'b0101;
	mem[3632] = 4'b0110;
	mem[3633] = 4'b0101;
	mem[3634] = 4'b0101;
	mem[3635] = 4'b0101;
	mem[3636] = 4'b0101;
	mem[3637] = 4'b0100;
	mem[3638] = 4'b0100;
	mem[3639] = 4'b0100;
	mem[3640] = 4'b0100;
	mem[3641] = 4'b0100;
	mem[3642] = 4'b0011;
	mem[3643] = 4'b0011;
	mem[3644] = 4'b0011;
	mem[3645] = 4'b0011;
	mem[3646] = 4'b0010;
	mem[3647] = 4'b0010;
	mem[3648] = 4'b0010;
	mem[3649] = 4'b0010;
	mem[3650] = 4'b0010;
	mem[3651] = 4'b0001;
	mem[3652] = 4'b0001;
	mem[3653] = 4'b0001;
	mem[3654] = 4'b0001;
	mem[3655] = 4'b0000;
	mem[3656] = 4'b0000;
	mem[3657] = 4'b0000;
	mem[3658] = 4'b0000;
	mem[3659] = 4'b1001;
	mem[3660] = 4'b1111;
	mem[3661] = 4'b1111;
	mem[3662] = 4'b1110;
	mem[3663] = 4'b1110;
	mem[3664] = 4'b1101;
	mem[3665] = 4'b1100;
	mem[3666] = 4'b1100;
	mem[3667] = 4'b1100;
	mem[3668] = 4'b1011;
	mem[3669] = 4'b1010;
	mem[3670] = 4'b1010;
	mem[3671] = 4'b1010;
	mem[3672] = 4'b1010;
	mem[3673] = 4'b1010;
	mem[3674] = 4'b1011;
	mem[3675] = 4'b1010;
	mem[3676] = 4'b1010;
	mem[3677] = 4'b1010;
	mem[3678] = 4'b1001;
	mem[3679] = 4'b1001;
	mem[3680] = 4'b1001;
	mem[3681] = 4'b1000;
	mem[3682] = 4'b1000;
	mem[3683] = 4'b1000;
	mem[3684] = 4'b1000;
	mem[3685] = 4'b0111;
	mem[3686] = 4'b0111;
	mem[3687] = 4'b0111;
	mem[3688] = 4'b0111;
	mem[3689] = 4'b0110;
	mem[3690] = 4'b0110;
	mem[3691] = 4'b0110;
	mem[3692] = 4'b0110;
	mem[3693] = 4'b0110;
	mem[3694] = 4'b0101;
	mem[3695] = 4'b0101;
	mem[3696] = 4'b0101;
	mem[3697] = 4'b0101;
	mem[3698] = 4'b0101;
	mem[3699] = 4'b0100;
	mem[3700] = 4'b0100;
	mem[3701] = 4'b0100;
	mem[3702] = 4'b0100;
	mem[3703] = 4'b0100;
	mem[3704] = 4'b0100;
	mem[3705] = 4'b0011;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b1001;
	mem[3716] = 4'b1111;
	mem[3717] = 4'b1111;
	mem[3718] = 4'b1111;
	mem[3719] = 4'b1111;
	mem[3720] = 4'b1110;
	mem[3721] = 4'b1110;
	mem[3722] = 4'b1110;
	mem[3723] = 4'b1110;
	mem[3724] = 4'b1101;
	mem[3725] = 4'b1101;
	mem[3726] = 4'b1101;
	mem[3727] = 4'b1101;
	mem[3728] = 4'b1101;
	mem[3729] = 4'b1100;
	mem[3730] = 4'b1100;
	mem[3731] = 4'b1100;
	mem[3732] = 4'b1100;
	mem[3733] = 4'b1011;
	mem[3734] = 4'b1011;
	mem[3735] = 4'b1011;
	mem[3736] = 4'b1011;
	mem[3737] = 4'b1010;
	mem[3738] = 4'b1001;
	mem[3739] = 4'b1001;
	mem[3740] = 4'b1001;
	mem[3741] = 4'b1001;
	mem[3742] = 4'b1010;
	mem[3743] = 4'b1010;
	mem[3744] = 4'b1001;
	mem[3745] = 4'b1001;
	mem[3746] = 4'b1001;
	mem[3747] = 4'b0111;
	mem[3748] = 4'b0111;
	mem[3749] = 4'b0111;
	mem[3750] = 4'b0111;
	mem[3751] = 4'b0111;
	mem[3752] = 4'b1000;
	mem[3753] = 4'b0111;
	mem[3754] = 4'b0111;
	mem[3755] = 4'b0111;
	mem[3756] = 4'b0111;
	mem[3757] = 4'b0110;
	mem[3758] = 4'b0110;
	mem[3759] = 4'b0111;
	mem[3760] = 4'b0110;
	mem[3761] = 4'b0101;
	mem[3762] = 4'b0101;
	mem[3763] = 4'b0101;
	mem[3764] = 4'b0101;
	mem[3765] = 4'b0100;
	mem[3766] = 4'b0100;
	mem[3767] = 4'b0100;
	mem[3768] = 4'b0100;
	mem[3769] = 4'b0100;
	mem[3770] = 4'b0011;
	mem[3771] = 4'b0011;
	mem[3772] = 4'b0011;
	mem[3773] = 4'b0011;
	mem[3774] = 4'b0010;
	mem[3775] = 4'b0010;
	mem[3776] = 4'b0010;
	mem[3777] = 4'b0010;
	mem[3778] = 4'b0010;
	mem[3779] = 4'b0001;
	mem[3780] = 4'b0001;
	mem[3781] = 4'b0001;
	mem[3782] = 4'b0001;
	mem[3783] = 4'b0000;
	mem[3784] = 4'b0000;
	mem[3785] = 4'b0000;
	mem[3786] = 4'b0000;
	mem[3787] = 4'b1001;
	mem[3788] = 4'b1111;
	mem[3789] = 4'b1111;
	mem[3790] = 4'b1110;
	mem[3791] = 4'b1110;
	mem[3792] = 4'b1110;
	mem[3793] = 4'b1011;
	mem[3794] = 4'b1011;
	mem[3795] = 4'b1011;
	mem[3796] = 4'b1011;
	mem[3797] = 4'b1011;
	mem[3798] = 4'b1100;
	mem[3799] = 4'b1100;
	mem[3800] = 4'b1010;
	mem[3801] = 4'b1010;
	mem[3802] = 4'b1011;
	mem[3803] = 4'b1010;
	mem[3804] = 4'b1010;
	mem[3805] = 4'b1010;
	mem[3806] = 4'b1001;
	mem[3807] = 4'b1001;
	mem[3808] = 4'b1001;
	mem[3809] = 4'b1001;
	mem[3810] = 4'b1000;
	mem[3811] = 4'b1000;
	mem[3812] = 4'b1000;
	mem[3813] = 4'b1000;
	mem[3814] = 4'b0111;
	mem[3815] = 4'b0111;
	mem[3816] = 4'b0111;
	mem[3817] = 4'b0111;
	mem[3818] = 4'b0110;
	mem[3819] = 4'b0110;
	mem[3820] = 4'b0110;
	mem[3821] = 4'b0110;
	mem[3822] = 4'b0110;
	mem[3823] = 4'b0101;
	mem[3824] = 4'b0101;
	mem[3825] = 4'b0101;
	mem[3826] = 4'b0101;
	mem[3827] = 4'b0101;
	mem[3828] = 4'b0100;
	mem[3829] = 4'b0100;
	mem[3830] = 4'b0100;
	mem[3831] = 4'b0100;
	mem[3832] = 4'b0100;
	mem[3833] = 4'b0011;
	mem[3834] = 4'b0000;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b1001;
	mem[3844] = 4'b1111;
	mem[3845] = 4'b1111;
	mem[3846] = 4'b1111;
	mem[3847] = 4'b1111;
	mem[3848] = 4'b1110;
	mem[3849] = 4'b1110;
	mem[3850] = 4'b1110;
	mem[3851] = 4'b1110;
	mem[3852] = 4'b1101;
	mem[3853] = 4'b1101;
	mem[3854] = 4'b1101;
	mem[3855] = 4'b1101;
	mem[3856] = 4'b1101;
	mem[3857] = 4'b1100;
	mem[3858] = 4'b1100;
	mem[3859] = 4'b1100;
	mem[3860] = 4'b1100;
	mem[3861] = 4'b1011;
	mem[3862] = 4'b1011;
	mem[3863] = 4'b1011;
	mem[3864] = 4'b1011;
	mem[3865] = 4'b1010;
	mem[3866] = 4'b1001;
	mem[3867] = 4'b1001;
	mem[3868] = 4'b1001;
	mem[3869] = 4'b1010;
	mem[3870] = 4'b1010;
	mem[3871] = 4'b1001;
	mem[3872] = 4'b1001;
	mem[3873] = 4'b1001;
	mem[3874] = 4'b1001;
	mem[3875] = 4'b1001;
	mem[3876] = 4'b0111;
	mem[3877] = 4'b0111;
	mem[3878] = 4'b0111;
	mem[3879] = 4'b0111;
	mem[3880] = 4'b0111;
	mem[3881] = 4'b0111;
	mem[3882] = 4'b0111;
	mem[3883] = 4'b0111;
	mem[3884] = 4'b0110;
	mem[3885] = 4'b0111;
	mem[3886] = 4'b0111;
	mem[3887] = 4'b0110;
	mem[3888] = 4'b0101;
	mem[3889] = 4'b0101;
	mem[3890] = 4'b0101;
	mem[3891] = 4'b0101;
	mem[3892] = 4'b0101;
	mem[3893] = 4'b0100;
	mem[3894] = 4'b0100;
	mem[3895] = 4'b0100;
	mem[3896] = 4'b0100;
	mem[3897] = 4'b0100;
	mem[3898] = 4'b0011;
	mem[3899] = 4'b0011;
	mem[3900] = 4'b0011;
	mem[3901] = 4'b0011;
	mem[3902] = 4'b0010;
	mem[3903] = 4'b0010;
	mem[3904] = 4'b0010;
	mem[3905] = 4'b0010;
	mem[3906] = 4'b0010;
	mem[3907] = 4'b0001;
	mem[3908] = 4'b0001;
	mem[3909] = 4'b0001;
	mem[3910] = 4'b0001;
	mem[3911] = 4'b0000;
	mem[3912] = 4'b0000;
	mem[3913] = 4'b0000;
	mem[3914] = 4'b0000;
	mem[3915] = 4'b1001;
	mem[3916] = 4'b1111;
	mem[3917] = 4'b1110;
	mem[3918] = 4'b1110;
	mem[3919] = 4'b1110;
	mem[3920] = 4'b1110;
	mem[3921] = 4'b1101;
	mem[3922] = 4'b1100;
	mem[3923] = 4'b1100;
	mem[3924] = 4'b1100;
	mem[3925] = 4'b1100;
	mem[3926] = 4'b1100;
	mem[3927] = 4'b1011;
	mem[3928] = 4'b1010;
	mem[3929] = 4'b1011;
	mem[3930] = 4'b1011;
	mem[3931] = 4'b1010;
	mem[3932] = 4'b1010;
	mem[3933] = 4'b1010;
	mem[3934] = 4'b1001;
	mem[3935] = 4'b1001;
	mem[3936] = 4'b1001;
	mem[3937] = 4'b1001;
	mem[3938] = 4'b1000;
	mem[3939] = 4'b1000;
	mem[3940] = 4'b1000;
	mem[3941] = 4'b1000;
	mem[3942] = 4'b0111;
	mem[3943] = 4'b0111;
	mem[3944] = 4'b0111;
	mem[3945] = 4'b0111;
	mem[3946] = 4'b0111;
	mem[3947] = 4'b0110;
	mem[3948] = 4'b0110;
	mem[3949] = 4'b0110;
	mem[3950] = 4'b0110;
	mem[3951] = 4'b0110;
	mem[3952] = 4'b0101;
	mem[3953] = 4'b0101;
	mem[3954] = 4'b0101;
	mem[3955] = 4'b0101;
	mem[3956] = 4'b0101;
	mem[3957] = 4'b0100;
	mem[3958] = 4'b0100;
	mem[3959] = 4'b0100;
	mem[3960] = 4'b0100;
	mem[3961] = 4'b0100;
	mem[3962] = 4'b0001;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b1001;
	mem[3972] = 4'b1111;
	mem[3973] = 4'b1111;
	mem[3974] = 4'b1111;
	mem[3975] = 4'b1111;
	mem[3976] = 4'b1110;
	mem[3977] = 4'b1110;
	mem[3978] = 4'b1110;
	mem[3979] = 4'b1110;
	mem[3980] = 4'b1101;
	mem[3981] = 4'b1101;
	mem[3982] = 4'b1101;
	mem[3983] = 4'b1101;
	mem[3984] = 4'b1101;
	mem[3985] = 4'b1100;
	mem[3986] = 4'b1100;
	mem[3987] = 4'b1100;
	mem[3988] = 4'b1100;
	mem[3989] = 4'b1011;
	mem[3990] = 4'b1011;
	mem[3991] = 4'b1011;
	mem[3992] = 4'b1011;
	mem[3993] = 4'b1010;
	mem[3994] = 4'b1001;
	mem[3995] = 4'b1001;
	mem[3996] = 4'b1001;
	mem[3997] = 4'b1010;
	mem[3998] = 4'b1001;
	mem[3999] = 4'b1001;
	mem[4000] = 4'b1001;
	mem[4001] = 4'b1001;
	mem[4002] = 4'b1001;
	mem[4003] = 4'b1000;
	mem[4004] = 4'b1000;
	mem[4005] = 4'b0111;
	mem[4006] = 4'b0111;
	mem[4007] = 4'b0111;
	mem[4008] = 4'b0111;
	mem[4009] = 4'b0111;
	mem[4010] = 4'b0111;
	mem[4011] = 4'b0111;
	mem[4012] = 4'b0110;
	mem[4013] = 4'b0110;
	mem[4014] = 4'b0110;
	mem[4015] = 4'b0110;
	mem[4016] = 4'b0101;
	mem[4017] = 4'b0101;
	mem[4018] = 4'b0101;
	mem[4019] = 4'b0101;
	mem[4020] = 4'b0101;
	mem[4021] = 4'b0100;
	mem[4022] = 4'b0100;
	mem[4023] = 4'b0100;
	mem[4024] = 4'b0100;
	mem[4025] = 4'b0100;
	mem[4026] = 4'b0011;
	mem[4027] = 4'b0011;
	mem[4028] = 4'b0011;
	mem[4029] = 4'b0011;
	mem[4030] = 4'b0010;
	mem[4031] = 4'b0010;
	mem[4032] = 4'b0010;
	mem[4033] = 4'b0010;
	mem[4034] = 4'b0010;
	mem[4035] = 4'b0001;
	mem[4036] = 4'b0001;
	mem[4037] = 4'b0001;
	mem[4038] = 4'b0001;
	mem[4039] = 4'b0000;
	mem[4040] = 4'b0000;
	mem[4041] = 4'b0000;
	mem[4042] = 4'b0000;
	mem[4043] = 4'b1001;
	mem[4044] = 4'b1110;
	mem[4045] = 4'b1101;
	mem[4046] = 4'b1101;
	mem[4047] = 4'b1101;
	mem[4048] = 4'b1110;
	mem[4049] = 4'b1101;
	mem[4050] = 4'b1101;
	mem[4051] = 4'b1101;
	mem[4052] = 4'b1100;
	mem[4053] = 4'b1011;
	mem[4054] = 4'b1011;
	mem[4055] = 4'b1010;
	mem[4056] = 4'b1010;
	mem[4057] = 4'b1011;
	mem[4058] = 4'b1011;
	mem[4059] = 4'b1010;
	mem[4060] = 4'b1010;
	mem[4061] = 4'b1010;
	mem[4062] = 4'b1010;
	mem[4063] = 4'b1001;
	mem[4064] = 4'b1001;
	mem[4065] = 4'b1001;
	mem[4066] = 4'b1001;
	mem[4067] = 4'b1000;
	mem[4068] = 4'b1000;
	mem[4069] = 4'b1000;
	mem[4070] = 4'b1000;
	mem[4071] = 4'b0111;
	mem[4072] = 4'b0111;
	mem[4073] = 4'b0111;
	mem[4074] = 4'b0111;
	mem[4075] = 4'b0111;
	mem[4076] = 4'b0110;
	mem[4077] = 4'b0110;
	mem[4078] = 4'b0110;
	mem[4079] = 4'b0110;
	mem[4080] = 4'b0110;
	mem[4081] = 4'b0101;
	mem[4082] = 4'b0101;
	mem[4083] = 4'b0101;
	mem[4084] = 4'b0101;
	mem[4085] = 4'b0101;
	mem[4086] = 4'b0101;
	mem[4087] = 4'b0100;
	mem[4088] = 4'b0100;
	mem[4089] = 4'b0100;
	mem[4090] = 4'b0001;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_3g (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0110;
	mem[4] = 4'b1001;
	mem[5] = 4'b1001;
	mem[6] = 4'b1001;
	mem[7] = 4'b1001;
	mem[8] = 4'b1001;
	mem[9] = 4'b1001;
	mem[10] = 4'b1001;
	mem[11] = 4'b1001;
	mem[12] = 4'b1001;
	mem[13] = 4'b1001;
	mem[14] = 4'b1001;
	mem[15] = 4'b1001;
	mem[16] = 4'b1001;
	mem[17] = 4'b1001;
	mem[18] = 4'b1001;
	mem[19] = 4'b1000;
	mem[20] = 4'b1001;
	mem[21] = 4'b1001;
	mem[22] = 4'b1001;
	mem[23] = 4'b1001;
	mem[24] = 4'b1000;
	mem[25] = 4'b1000;
	mem[26] = 4'b1000;
	mem[27] = 4'b1000;
	mem[28] = 4'b1000;
	mem[29] = 4'b1001;
	mem[30] = 4'b1000;
	mem[31] = 4'b1000;
	mem[32] = 4'b1000;
	mem[33] = 4'b1000;
	mem[34] = 4'b1000;
	mem[35] = 4'b1000;
	mem[36] = 4'b1000;
	mem[37] = 4'b1000;
	mem[38] = 4'b0111;
	mem[39] = 4'b0111;
	mem[40] = 4'b0111;
	mem[41] = 4'b1000;
	mem[42] = 4'b1000;
	mem[43] = 4'b1000;
	mem[44] = 4'b1000;
	mem[45] = 4'b1000;
	mem[46] = 4'b1000;
	mem[47] = 4'b1000;
	mem[48] = 4'b1000;
	mem[49] = 4'b1000;
	mem[50] = 4'b1000;
	mem[51] = 4'b1000;
	mem[52] = 4'b0111;
	mem[53] = 4'b1000;
	mem[54] = 4'b1000;
	mem[55] = 4'b1000;
	mem[56] = 4'b1000;
	mem[57] = 4'b0111;
	mem[58] = 4'b0111;
	mem[59] = 4'b0111;
	mem[60] = 4'b0111;
	mem[61] = 4'b0111;
	mem[62] = 4'b0111;
	mem[63] = 4'b0111;
	mem[64] = 4'b0111;
	mem[65] = 4'b0111;
	mem[66] = 4'b0111;
	mem[67] = 4'b0111;
	mem[68] = 4'b0111;
	mem[69] = 4'b0110;
	mem[70] = 4'b0011;
	mem[71] = 4'b0000;
	mem[72] = 4'b0000;
	mem[73] = 4'b0000;
	mem[74] = 4'b0000;
	mem[75] = 4'b0101;
	mem[76] = 4'b1000;
	mem[77] = 4'b1000;
	mem[78] = 4'b1000;
	mem[79] = 4'b1000;
	mem[80] = 4'b1000;
	mem[81] = 4'b1000;
	mem[82] = 4'b1000;
	mem[83] = 4'b1000;
	mem[84] = 4'b0111;
	mem[85] = 4'b0111;
	mem[86] = 4'b0111;
	mem[87] = 4'b1000;
	mem[88] = 4'b1000;
	mem[89] = 4'b0111;
	mem[90] = 4'b0111;
	mem[91] = 4'b0111;
	mem[92] = 4'b0111;
	mem[93] = 4'b0111;
	mem[94] = 4'b0111;
	mem[95] = 4'b0110;
	mem[96] = 4'b0110;
	mem[97] = 4'b0110;
	mem[98] = 4'b0110;
	mem[99] = 4'b0110;
	mem[100] = 4'b0110;
	mem[101] = 4'b0110;
	mem[102] = 4'b0110;
	mem[103] = 4'b0110;
	mem[104] = 4'b0101;
	mem[105] = 4'b0101;
	mem[106] = 4'b0101;
	mem[107] = 4'b0101;
	mem[108] = 4'b0101;
	mem[109] = 4'b0101;
	mem[110] = 4'b0101;
	mem[111] = 4'b0101;
	mem[112] = 4'b0101;
	mem[113] = 4'b0101;
	mem[114] = 4'b0101;
	mem[115] = 4'b0101;
	mem[116] = 4'b0101;
	mem[117] = 4'b0101;
	mem[118] = 4'b0101;
	mem[119] = 4'b0100;
	mem[120] = 4'b0100;
	mem[121] = 4'b0100;
	mem[122] = 4'b0001;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b0000;
	mem[132] = 4'b0000;
	mem[133] = 4'b0000;
	mem[134] = 4'b0000;
	mem[135] = 4'b0000;
	mem[136] = 4'b0000;
	mem[137] = 4'b0001;
	mem[138] = 4'b0001;
	mem[139] = 4'b0001;
	mem[140] = 4'b0001;
	mem[141] = 4'b0001;
	mem[142] = 4'b0010;
	mem[143] = 4'b0011;
	mem[144] = 4'b0011;
	mem[145] = 4'b0011;
	mem[146] = 4'b0011;
	mem[147] = 4'b0011;
	mem[148] = 4'b0100;
	mem[149] = 4'b0100;
	mem[150] = 4'b0100;
	mem[151] = 4'b0100;
	mem[152] = 4'b0100;
	mem[153] = 4'b0101;
	mem[154] = 4'b0101;
	mem[155] = 4'b0101;
	mem[156] = 4'b0110;
	mem[157] = 4'b0110;
	mem[158] = 4'b0110;
	mem[159] = 4'b0111;
	mem[160] = 4'b1000;
	mem[161] = 4'b1000;
	mem[162] = 4'b1000;
	mem[163] = 4'b1000;
	mem[164] = 4'b1000;
	mem[165] = 4'b1001;
	mem[166] = 4'b1000;
	mem[167] = 4'b1000;
	mem[168] = 4'b1000;
	mem[169] = 4'b1001;
	mem[170] = 4'b1010;
	mem[171] = 4'b1011;
	mem[172] = 4'b1011;
	mem[173] = 4'b1011;
	mem[174] = 4'b1011;
	mem[175] = 4'b1011;
	mem[176] = 4'b1100;
	mem[177] = 4'b1100;
	mem[178] = 4'b1100;
	mem[179] = 4'b1100;
	mem[180] = 4'b1100;
	mem[181] = 4'b1101;
	mem[182] = 4'b1110;
	mem[183] = 4'b1110;
	mem[184] = 4'b1110;
	mem[185] = 4'b1110;
	mem[186] = 4'b1110;
	mem[187] = 4'b1111;
	mem[188] = 4'b1111;
	mem[189] = 4'b1111;
	mem[190] = 4'b1111;
	mem[191] = 4'b1111;
	mem[192] = 4'b1111;
	mem[193] = 4'b1111;
	mem[194] = 4'b1111;
	mem[195] = 4'b1111;
	mem[196] = 4'b1111;
	mem[197] = 4'b1111;
	mem[198] = 4'b0110;
	mem[199] = 4'b0000;
	mem[200] = 4'b0000;
	mem[201] = 4'b0000;
	mem[202] = 4'b0000;
	mem[203] = 4'b0000;
	mem[204] = 4'b0001;
	mem[205] = 4'b0001;
	mem[206] = 4'b0001;
	mem[207] = 4'b0000;
	mem[208] = 4'b0000;
	mem[209] = 4'b0001;
	mem[210] = 4'b0001;
	mem[211] = 4'b0000;
	mem[212] = 4'b0001;
	mem[213] = 4'b0010;
	mem[214] = 4'b0010;
	mem[215] = 4'b0010;
	mem[216] = 4'b0001;
	mem[217] = 4'b0001;
	mem[218] = 4'b0001;
	mem[219] = 4'b0001;
	mem[220] = 4'b0001;
	mem[221] = 4'b0001;
	mem[222] = 4'b0010;
	mem[223] = 4'b0010;
	mem[224] = 4'b0010;
	mem[225] = 4'b0010;
	mem[226] = 4'b0010;
	mem[227] = 4'b0010;
	mem[228] = 4'b0010;
	mem[229] = 4'b0010;
	mem[230] = 4'b0010;
	mem[231] = 4'b0011;
	mem[232] = 4'b0011;
	mem[233] = 4'b0011;
	mem[234] = 4'b0011;
	mem[235] = 4'b0011;
	mem[236] = 4'b0011;
	mem[237] = 4'b0011;
	mem[238] = 4'b0011;
	mem[239] = 4'b0011;
	mem[240] = 4'b0100;
	mem[241] = 4'b0100;
	mem[242] = 4'b0100;
	mem[243] = 4'b0100;
	mem[244] = 4'b0100;
	mem[245] = 4'b0100;
	mem[246] = 4'b0100;
	mem[247] = 4'b0100;
	mem[248] = 4'b0100;
	mem[249] = 4'b0100;
	mem[250] = 4'b0001;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0000;
	mem[260] = 4'b0000;
	mem[261] = 4'b0000;
	mem[262] = 4'b0000;
	mem[263] = 4'b0000;
	mem[264] = 4'b0000;
	mem[265] = 4'b0001;
	mem[266] = 4'b0001;
	mem[267] = 4'b0001;
	mem[268] = 4'b0001;
	mem[269] = 4'b0001;
	mem[270] = 4'b0010;
	mem[271] = 4'b0011;
	mem[272] = 4'b0011;
	mem[273] = 4'b0011;
	mem[274] = 4'b0011;
	mem[275] = 4'b0011;
	mem[276] = 4'b0100;
	mem[277] = 4'b0100;
	mem[278] = 4'b0100;
	mem[279] = 4'b0100;
	mem[280] = 4'b0100;
	mem[281] = 4'b0101;
	mem[282] = 4'b0101;
	mem[283] = 4'b0101;
	mem[284] = 4'b0101;
	mem[285] = 4'b0110;
	mem[286] = 4'b0110;
	mem[287] = 4'b0111;
	mem[288] = 4'b1000;
	mem[289] = 4'b1000;
	mem[290] = 4'b1000;
	mem[291] = 4'b1000;
	mem[292] = 4'b1000;
	mem[293] = 4'b1000;
	mem[294] = 4'b1000;
	mem[295] = 4'b1000;
	mem[296] = 4'b1001;
	mem[297] = 4'b1001;
	mem[298] = 4'b1010;
	mem[299] = 4'b1011;
	mem[300] = 4'b1011;
	mem[301] = 4'b1011;
	mem[302] = 4'b1011;
	mem[303] = 4'b1011;
	mem[304] = 4'b1100;
	mem[305] = 4'b1100;
	mem[306] = 4'b1100;
	mem[307] = 4'b1100;
	mem[308] = 4'b1100;
	mem[309] = 4'b1101;
	mem[310] = 4'b1110;
	mem[311] = 4'b1110;
	mem[312] = 4'b1110;
	mem[313] = 4'b1110;
	mem[314] = 4'b1110;
	mem[315] = 4'b1111;
	mem[316] = 4'b1111;
	mem[317] = 4'b1111;
	mem[318] = 4'b1111;
	mem[319] = 4'b1111;
	mem[320] = 4'b1111;
	mem[321] = 4'b1111;
	mem[322] = 4'b1111;
	mem[323] = 4'b1111;
	mem[324] = 4'b1111;
	mem[325] = 4'b1111;
	mem[326] = 4'b0110;
	mem[327] = 4'b0000;
	mem[328] = 4'b0000;
	mem[329] = 4'b0000;
	mem[330] = 4'b0000;
	mem[331] = 4'b0000;
	mem[332] = 4'b0001;
	mem[333] = 4'b0000;
	mem[334] = 4'b0000;
	mem[335] = 4'b0001;
	mem[336] = 4'b0001;
	mem[337] = 4'b0001;
	mem[338] = 4'b0001;
	mem[339] = 4'b0001;
	mem[340] = 4'b0001;
	mem[341] = 4'b0001;
	mem[342] = 4'b0001;
	mem[343] = 4'b0001;
	mem[344] = 4'b0001;
	mem[345] = 4'b0001;
	mem[346] = 4'b0001;
	mem[347] = 4'b0010;
	mem[348] = 4'b0010;
	mem[349] = 4'b0010;
	mem[350] = 4'b0010;
	mem[351] = 4'b0010;
	mem[352] = 4'b0010;
	mem[353] = 4'b0010;
	mem[354] = 4'b0010;
	mem[355] = 4'b0010;
	mem[356] = 4'b0011;
	mem[357] = 4'b0011;
	mem[358] = 4'b0011;
	mem[359] = 4'b0011;
	mem[360] = 4'b0011;
	mem[361] = 4'b0011;
	mem[362] = 4'b0011;
	mem[363] = 4'b0011;
	mem[364] = 4'b0011;
	mem[365] = 4'b0011;
	mem[366] = 4'b0100;
	mem[367] = 4'b0100;
	mem[368] = 4'b0100;
	mem[369] = 4'b0100;
	mem[370] = 4'b0100;
	mem[371] = 4'b0100;
	mem[372] = 4'b0100;
	mem[373] = 4'b0100;
	mem[374] = 4'b0100;
	mem[375] = 4'b0101;
	mem[376] = 4'b0101;
	mem[377] = 4'b0101;
	mem[378] = 4'b0001;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0000;
	mem[388] = 4'b0000;
	mem[389] = 4'b0000;
	mem[390] = 4'b0000;
	mem[391] = 4'b0000;
	mem[392] = 4'b0000;
	mem[393] = 4'b0001;
	mem[394] = 4'b0001;
	mem[395] = 4'b0001;
	mem[396] = 4'b0001;
	mem[397] = 4'b0001;
	mem[398] = 4'b0010;
	mem[399] = 4'b0011;
	mem[400] = 4'b0011;
	mem[401] = 4'b0011;
	mem[402] = 4'b0011;
	mem[403] = 4'b0011;
	mem[404] = 4'b0100;
	mem[405] = 4'b0100;
	mem[406] = 4'b0100;
	mem[407] = 4'b0100;
	mem[408] = 4'b0100;
	mem[409] = 4'b0101;
	mem[410] = 4'b0101;
	mem[411] = 4'b0101;
	mem[412] = 4'b0101;
	mem[413] = 4'b0101;
	mem[414] = 4'b0110;
	mem[415] = 4'b0111;
	mem[416] = 4'b1000;
	mem[417] = 4'b1000;
	mem[418] = 4'b1000;
	mem[419] = 4'b1000;
	mem[420] = 4'b1000;
	mem[421] = 4'b1000;
	mem[422] = 4'b1000;
	mem[423] = 4'b1000;
	mem[424] = 4'b1001;
	mem[425] = 4'b1001;
	mem[426] = 4'b1010;
	mem[427] = 4'b1011;
	mem[428] = 4'b1011;
	mem[429] = 4'b1011;
	mem[430] = 4'b1011;
	mem[431] = 4'b1011;
	mem[432] = 4'b1100;
	mem[433] = 4'b1100;
	mem[434] = 4'b1100;
	mem[435] = 4'b1100;
	mem[436] = 4'b1100;
	mem[437] = 4'b1101;
	mem[438] = 4'b1110;
	mem[439] = 4'b1110;
	mem[440] = 4'b1110;
	mem[441] = 4'b1110;
	mem[442] = 4'b1110;
	mem[443] = 4'b1111;
	mem[444] = 4'b1111;
	mem[445] = 4'b1111;
	mem[446] = 4'b1111;
	mem[447] = 4'b1111;
	mem[448] = 4'b1111;
	mem[449] = 4'b1111;
	mem[450] = 4'b1111;
	mem[451] = 4'b1111;
	mem[452] = 4'b1111;
	mem[453] = 4'b1111;
	mem[454] = 4'b0110;
	mem[455] = 4'b0000;
	mem[456] = 4'b0000;
	mem[457] = 4'b0000;
	mem[458] = 4'b0000;
	mem[459] = 4'b0001;
	mem[460] = 4'b0001;
	mem[461] = 4'b0000;
	mem[462] = 4'b0000;
	mem[463] = 4'b0001;
	mem[464] = 4'b0001;
	mem[465] = 4'b0001;
	mem[466] = 4'b0001;
	mem[467] = 4'b0010;
	mem[468] = 4'b0001;
	mem[469] = 4'b0001;
	mem[470] = 4'b0001;
	mem[471] = 4'b0001;
	mem[472] = 4'b0001;
	mem[473] = 4'b0010;
	mem[474] = 4'b0010;
	mem[475] = 4'b0010;
	mem[476] = 4'b0010;
	mem[477] = 4'b0010;
	mem[478] = 4'b0010;
	mem[479] = 4'b0010;
	mem[480] = 4'b0010;
	mem[481] = 4'b0010;
	mem[482] = 4'b0011;
	mem[483] = 4'b0011;
	mem[484] = 4'b0011;
	mem[485] = 4'b0011;
	mem[486] = 4'b0011;
	mem[487] = 4'b0011;
	mem[488] = 4'b0011;
	mem[489] = 4'b0011;
	mem[490] = 4'b0011;
	mem[491] = 4'b0100;
	mem[492] = 4'b0100;
	mem[493] = 4'b0100;
	mem[494] = 4'b0100;
	mem[495] = 4'b0100;
	mem[496] = 4'b0100;
	mem[497] = 4'b0100;
	mem[498] = 4'b0100;
	mem[499] = 4'b0100;
	mem[500] = 4'b0101;
	mem[501] = 4'b0101;
	mem[502] = 4'b0101;
	mem[503] = 4'b0101;
	mem[504] = 4'b0101;
	mem[505] = 4'b0101;
	mem[506] = 4'b0001;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0000;
	mem[516] = 4'b0000;
	mem[517] = 4'b0000;
	mem[518] = 4'b0000;
	mem[519] = 4'b0000;
	mem[520] = 4'b0000;
	mem[521] = 4'b0001;
	mem[522] = 4'b0001;
	mem[523] = 4'b0001;
	mem[524] = 4'b0001;
	mem[525] = 4'b0001;
	mem[526] = 4'b0010;
	mem[527] = 4'b0011;
	mem[528] = 4'b0011;
	mem[529] = 4'b0011;
	mem[530] = 4'b0011;
	mem[531] = 4'b0011;
	mem[532] = 4'b0100;
	mem[533] = 4'b0100;
	mem[534] = 4'b0100;
	mem[535] = 4'b0100;
	mem[536] = 4'b0100;
	mem[537] = 4'b0101;
	mem[538] = 4'b0110;
	mem[539] = 4'b0101;
	mem[540] = 4'b0101;
	mem[541] = 4'b0101;
	mem[542] = 4'b0101;
	mem[543] = 4'b0111;
	mem[544] = 4'b1000;
	mem[545] = 4'b1000;
	mem[546] = 4'b0111;
	mem[547] = 4'b0111;
	mem[548] = 4'b0111;
	mem[549] = 4'b1000;
	mem[550] = 4'b1000;
	mem[551] = 4'b1000;
	mem[552] = 4'b1010;
	mem[553] = 4'b1001;
	mem[554] = 4'b1010;
	mem[555] = 4'b1011;
	mem[556] = 4'b1011;
	mem[557] = 4'b1011;
	mem[558] = 4'b1011;
	mem[559] = 4'b1011;
	mem[560] = 4'b1100;
	mem[561] = 4'b1100;
	mem[562] = 4'b1100;
	mem[563] = 4'b1100;
	mem[564] = 4'b1100;
	mem[565] = 4'b1101;
	mem[566] = 4'b1110;
	mem[567] = 4'b1110;
	mem[568] = 4'b1110;
	mem[569] = 4'b1110;
	mem[570] = 4'b1110;
	mem[571] = 4'b1111;
	mem[572] = 4'b1111;
	mem[573] = 4'b1111;
	mem[574] = 4'b1111;
	mem[575] = 4'b1111;
	mem[576] = 4'b1111;
	mem[577] = 4'b1111;
	mem[578] = 4'b1111;
	mem[579] = 4'b1111;
	mem[580] = 4'b1111;
	mem[581] = 4'b1111;
	mem[582] = 4'b0110;
	mem[583] = 4'b0000;
	mem[584] = 4'b0000;
	mem[585] = 4'b0001;
	mem[586] = 4'b0001;
	mem[587] = 4'b0001;
	mem[588] = 4'b0001;
	mem[589] = 4'b0001;
	mem[590] = 4'b0001;
	mem[591] = 4'b0001;
	mem[592] = 4'b0001;
	mem[593] = 4'b0010;
	mem[594] = 4'b0001;
	mem[595] = 4'b0010;
	mem[596] = 4'b0010;
	mem[597] = 4'b0001;
	mem[598] = 4'b0010;
	mem[599] = 4'b0010;
	mem[600] = 4'b0010;
	mem[601] = 4'b0010;
	mem[602] = 4'b0010;
	mem[603] = 4'b0010;
	mem[604] = 4'b0010;
	mem[605] = 4'b0010;
	mem[606] = 4'b0010;
	mem[607] = 4'b0011;
	mem[608] = 4'b0011;
	mem[609] = 4'b0011;
	mem[610] = 4'b0011;
	mem[611] = 4'b0011;
	mem[612] = 4'b0011;
	mem[613] = 4'b0011;
	mem[614] = 4'b0011;
	mem[615] = 4'b0011;
	mem[616] = 4'b0100;
	mem[617] = 4'b0100;
	mem[618] = 4'b0100;
	mem[619] = 4'b0100;
	mem[620] = 4'b0100;
	mem[621] = 4'b0100;
	mem[622] = 4'b0100;
	mem[623] = 4'b0100;
	mem[624] = 4'b0100;
	mem[625] = 4'b0100;
	mem[626] = 4'b0101;
	mem[627] = 4'b0101;
	mem[628] = 4'b0101;
	mem[629] = 4'b0101;
	mem[630] = 4'b0101;
	mem[631] = 4'b0101;
	mem[632] = 4'b0101;
	mem[633] = 4'b0101;
	mem[634] = 4'b0001;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0000;
	mem[644] = 4'b0000;
	mem[645] = 4'b0000;
	mem[646] = 4'b0000;
	mem[647] = 4'b0000;
	mem[648] = 4'b0000;
	mem[649] = 4'b0001;
	mem[650] = 4'b0001;
	mem[651] = 4'b0001;
	mem[652] = 4'b0001;
	mem[653] = 4'b0001;
	mem[654] = 4'b0010;
	mem[655] = 4'b0011;
	mem[656] = 4'b0011;
	mem[657] = 4'b0011;
	mem[658] = 4'b0011;
	mem[659] = 4'b0011;
	mem[660] = 4'b0100;
	mem[661] = 4'b0100;
	mem[662] = 4'b0100;
	mem[663] = 4'b0101;
	mem[664] = 4'b0100;
	mem[665] = 4'b0101;
	mem[666] = 4'b0110;
	mem[667] = 4'b0101;
	mem[668] = 4'b0101;
	mem[669] = 4'b0101;
	mem[670] = 4'b0101;
	mem[671] = 4'b0110;
	mem[672] = 4'b0111;
	mem[673] = 4'b0111;
	mem[674] = 4'b0111;
	mem[675] = 4'b0111;
	mem[676] = 4'b0111;
	mem[677] = 4'b1000;
	mem[678] = 4'b1000;
	mem[679] = 4'b1001;
	mem[680] = 4'b1001;
	mem[681] = 4'b1001;
	mem[682] = 4'b1010;
	mem[683] = 4'b1011;
	mem[684] = 4'b1011;
	mem[685] = 4'b1011;
	mem[686] = 4'b1011;
	mem[687] = 4'b1011;
	mem[688] = 4'b1100;
	mem[689] = 4'b1100;
	mem[690] = 4'b1100;
	mem[691] = 4'b1100;
	mem[692] = 4'b1100;
	mem[693] = 4'b1101;
	mem[694] = 4'b1110;
	mem[695] = 4'b1110;
	mem[696] = 4'b1110;
	mem[697] = 4'b1110;
	mem[698] = 4'b1110;
	mem[699] = 4'b1111;
	mem[700] = 4'b1111;
	mem[701] = 4'b1111;
	mem[702] = 4'b1111;
	mem[703] = 4'b1111;
	mem[704] = 4'b1111;
	mem[705] = 4'b1111;
	mem[706] = 4'b1111;
	mem[707] = 4'b1111;
	mem[708] = 4'b1111;
	mem[709] = 4'b1111;
	mem[710] = 4'b0110;
	mem[711] = 4'b0000;
	mem[712] = 4'b0000;
	mem[713] = 4'b0000;
	mem[714] = 4'b0001;
	mem[715] = 4'b0001;
	mem[716] = 4'b0001;
	mem[717] = 4'b0010;
	mem[718] = 4'b0001;
	mem[719] = 4'b0001;
	mem[720] = 4'b0001;
	mem[721] = 4'b0001;
	mem[722] = 4'b0010;
	mem[723] = 4'b0011;
	mem[724] = 4'b0010;
	mem[725] = 4'b0010;
	mem[726] = 4'b0010;
	mem[727] = 4'b0010;
	mem[728] = 4'b0010;
	mem[729] = 4'b0010;
	mem[730] = 4'b0010;
	mem[731] = 4'b0010;
	mem[732] = 4'b0010;
	mem[733] = 4'b0011;
	mem[734] = 4'b0011;
	mem[735] = 4'b0011;
	mem[736] = 4'b0011;
	mem[737] = 4'b0011;
	mem[738] = 4'b0011;
	mem[739] = 4'b0011;
	mem[740] = 4'b0011;
	mem[741] = 4'b0011;
	mem[742] = 4'b0100;
	mem[743] = 4'b0100;
	mem[744] = 4'b0100;
	mem[745] = 4'b0100;
	mem[746] = 4'b0100;
	mem[747] = 4'b0100;
	mem[748] = 4'b0100;
	mem[749] = 4'b0100;
	mem[750] = 4'b0100;
	mem[751] = 4'b0101;
	mem[752] = 4'b0101;
	mem[753] = 4'b0101;
	mem[754] = 4'b0101;
	mem[755] = 4'b0101;
	mem[756] = 4'b0101;
	mem[757] = 4'b0101;
	mem[758] = 4'b0101;
	mem[759] = 4'b0101;
	mem[760] = 4'b0110;
	mem[761] = 4'b0101;
	mem[762] = 4'b0001;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0000;
	mem[772] = 4'b0000;
	mem[773] = 4'b0000;
	mem[774] = 4'b0000;
	mem[775] = 4'b0000;
	mem[776] = 4'b0000;
	mem[777] = 4'b0001;
	mem[778] = 4'b0001;
	mem[779] = 4'b0001;
	mem[780] = 4'b0001;
	mem[781] = 4'b0001;
	mem[782] = 4'b0010;
	mem[783] = 4'b0011;
	mem[784] = 4'b0011;
	mem[785] = 4'b0011;
	mem[786] = 4'b0011;
	mem[787] = 4'b0011;
	mem[788] = 4'b0100;
	mem[789] = 4'b0100;
	mem[790] = 4'b0100;
	mem[791] = 4'b0101;
	mem[792] = 4'b0101;
	mem[793] = 4'b0101;
	mem[794] = 4'b0110;
	mem[795] = 4'b0110;
	mem[796] = 4'b0101;
	mem[797] = 4'b0101;
	mem[798] = 4'b0101;
	mem[799] = 4'b0110;
	mem[800] = 4'b0111;
	mem[801] = 4'b0111;
	mem[802] = 4'b0111;
	mem[803] = 4'b0111;
	mem[804] = 4'b0111;
	mem[805] = 4'b1000;
	mem[806] = 4'b1001;
	mem[807] = 4'b1010;
	mem[808] = 4'b1001;
	mem[809] = 4'b1001;
	mem[810] = 4'b1010;
	mem[811] = 4'b1011;
	mem[812] = 4'b1011;
	mem[813] = 4'b1011;
	mem[814] = 4'b1011;
	mem[815] = 4'b1011;
	mem[816] = 4'b1100;
	mem[817] = 4'b1100;
	mem[818] = 4'b1100;
	mem[819] = 4'b1100;
	mem[820] = 4'b1100;
	mem[821] = 4'b1101;
	mem[822] = 4'b1110;
	mem[823] = 4'b1110;
	mem[824] = 4'b1110;
	mem[825] = 4'b1110;
	mem[826] = 4'b1110;
	mem[827] = 4'b1111;
	mem[828] = 4'b1111;
	mem[829] = 4'b1111;
	mem[830] = 4'b1111;
	mem[831] = 4'b1111;
	mem[832] = 4'b1111;
	mem[833] = 4'b1111;
	mem[834] = 4'b1111;
	mem[835] = 4'b1111;
	mem[836] = 4'b1111;
	mem[837] = 4'b1110;
	mem[838] = 4'b0110;
	mem[839] = 4'b0001;
	mem[840] = 4'b0001;
	mem[841] = 4'b0001;
	mem[842] = 4'b0001;
	mem[843] = 4'b0010;
	mem[844] = 4'b0001;
	mem[845] = 4'b0001;
	mem[846] = 4'b0010;
	mem[847] = 4'b0010;
	mem[848] = 4'b0001;
	mem[849] = 4'b0010;
	mem[850] = 4'b0010;
	mem[851] = 4'b0010;
	mem[852] = 4'b0010;
	mem[853] = 4'b0010;
	mem[854] = 4'b0010;
	mem[855] = 4'b0010;
	mem[856] = 4'b0010;
	mem[857] = 4'b0010;
	mem[858] = 4'b0011;
	mem[859] = 4'b0011;
	mem[860] = 4'b0011;
	mem[861] = 4'b0011;
	mem[862] = 4'b0011;
	mem[863] = 4'b0011;
	mem[864] = 4'b0011;
	mem[865] = 4'b0011;
	mem[866] = 4'b0011;
	mem[867] = 4'b0100;
	mem[868] = 4'b0100;
	mem[869] = 4'b0100;
	mem[870] = 4'b0100;
	mem[871] = 4'b0100;
	mem[872] = 4'b0100;
	mem[873] = 4'b0100;
	mem[874] = 4'b0100;
	mem[875] = 4'b0100;
	mem[876] = 4'b0101;
	mem[877] = 4'b0101;
	mem[878] = 4'b0101;
	mem[879] = 4'b0101;
	mem[880] = 4'b0101;
	mem[881] = 4'b0101;
	mem[882] = 4'b0101;
	mem[883] = 4'b0101;
	mem[884] = 4'b0101;
	mem[885] = 4'b0101;
	mem[886] = 4'b0110;
	mem[887] = 4'b0110;
	mem[888] = 4'b0110;
	mem[889] = 4'b0110;
	mem[890] = 4'b0001;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0000;
	mem[900] = 4'b0000;
	mem[901] = 4'b0000;
	mem[902] = 4'b0000;
	mem[903] = 4'b0000;
	mem[904] = 4'b0000;
	mem[905] = 4'b0001;
	mem[906] = 4'b0001;
	mem[907] = 4'b0001;
	mem[908] = 4'b0001;
	mem[909] = 4'b0001;
	mem[910] = 4'b0010;
	mem[911] = 4'b0011;
	mem[912] = 4'b0011;
	mem[913] = 4'b0011;
	mem[914] = 4'b0011;
	mem[915] = 4'b0011;
	mem[916] = 4'b0100;
	mem[917] = 4'b0100;
	mem[918] = 4'b0101;
	mem[919] = 4'b0101;
	mem[920] = 4'b0100;
	mem[921] = 4'b0101;
	mem[922] = 4'b0110;
	mem[923] = 4'b0110;
	mem[924] = 4'b0110;
	mem[925] = 4'b0110;
	mem[926] = 4'b0101;
	mem[927] = 4'b0110;
	mem[928] = 4'b0111;
	mem[929] = 4'b0111;
	mem[930] = 4'b0111;
	mem[931] = 4'b0111;
	mem[932] = 4'b0111;
	mem[933] = 4'b1001;
	mem[934] = 4'b1010;
	mem[935] = 4'b1001;
	mem[936] = 4'b1001;
	mem[937] = 4'b1001;
	mem[938] = 4'b1010;
	mem[939] = 4'b1011;
	mem[940] = 4'b1011;
	mem[941] = 4'b1011;
	mem[942] = 4'b1011;
	mem[943] = 4'b1011;
	mem[944] = 4'b1100;
	mem[945] = 4'b1100;
	mem[946] = 4'b1100;
	mem[947] = 4'b1100;
	mem[948] = 4'b1100;
	mem[949] = 4'b1101;
	mem[950] = 4'b1110;
	mem[951] = 4'b1110;
	mem[952] = 4'b1110;
	mem[953] = 4'b1110;
	mem[954] = 4'b1110;
	mem[955] = 4'b1111;
	mem[956] = 4'b1111;
	mem[957] = 4'b1111;
	mem[958] = 4'b1111;
	mem[959] = 4'b1111;
	mem[960] = 4'b1111;
	mem[961] = 4'b1111;
	mem[962] = 4'b1111;
	mem[963] = 4'b1111;
	mem[964] = 4'b1110;
	mem[965] = 4'b1101;
	mem[966] = 4'b0110;
	mem[967] = 4'b0001;
	mem[968] = 4'b0001;
	mem[969] = 4'b0001;
	mem[970] = 4'b0010;
	mem[971] = 4'b0001;
	mem[972] = 4'b0010;
	mem[973] = 4'b0010;
	mem[974] = 4'b0010;
	mem[975] = 4'b0010;
	mem[976] = 4'b0010;
	mem[977] = 4'b0010;
	mem[978] = 4'b0010;
	mem[979] = 4'b0010;
	mem[980] = 4'b0010;
	mem[981] = 4'b0010;
	mem[982] = 4'b0010;
	mem[983] = 4'b0010;
	mem[984] = 4'b0011;
	mem[985] = 4'b0011;
	mem[986] = 4'b0011;
	mem[987] = 4'b0011;
	mem[988] = 4'b0011;
	mem[989] = 4'b0011;
	mem[990] = 4'b0011;
	mem[991] = 4'b0011;
	mem[992] = 4'b0011;
	mem[993] = 4'b0100;
	mem[994] = 4'b0100;
	mem[995] = 4'b0100;
	mem[996] = 4'b0100;
	mem[997] = 4'b0100;
	mem[998] = 4'b0100;
	mem[999] = 4'b0100;
	mem[1000] = 4'b0100;
	mem[1001] = 4'b0100;
	mem[1002] = 4'b0101;
	mem[1003] = 4'b0101;
	mem[1004] = 4'b0101;
	mem[1005] = 4'b0101;
	mem[1006] = 4'b0101;
	mem[1007] = 4'b0101;
	mem[1008] = 4'b0101;
	mem[1009] = 4'b0101;
	mem[1010] = 4'b0101;
	mem[1011] = 4'b0110;
	mem[1012] = 4'b0110;
	mem[1013] = 4'b0110;
	mem[1014] = 4'b0110;
	mem[1015] = 4'b0110;
	mem[1016] = 4'b0110;
	mem[1017] = 4'b0110;
	mem[1018] = 4'b0001;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0000;
	mem[1028] = 4'b0000;
	mem[1029] = 4'b0000;
	mem[1030] = 4'b0000;
	mem[1031] = 4'b0000;
	mem[1032] = 4'b0000;
	mem[1033] = 4'b0001;
	mem[1034] = 4'b0001;
	mem[1035] = 4'b0001;
	mem[1036] = 4'b0001;
	mem[1037] = 4'b0001;
	mem[1038] = 4'b0010;
	mem[1039] = 4'b0011;
	mem[1040] = 4'b0011;
	mem[1041] = 4'b0011;
	mem[1042] = 4'b0011;
	mem[1043] = 4'b0100;
	mem[1044] = 4'b0101;
	mem[1045] = 4'b0101;
	mem[1046] = 4'b0101;
	mem[1047] = 4'b0100;
	mem[1048] = 4'b0100;
	mem[1049] = 4'b0101;
	mem[1050] = 4'b0110;
	mem[1051] = 4'b0110;
	mem[1052] = 4'b0110;
	mem[1053] = 4'b0110;
	mem[1054] = 4'b0110;
	mem[1055] = 4'b0111;
	mem[1056] = 4'b0111;
	mem[1057] = 4'b0111;
	mem[1058] = 4'b0111;
	mem[1059] = 4'b1000;
	mem[1060] = 4'b1000;
	mem[1061] = 4'b1001;
	mem[1062] = 4'b1001;
	mem[1063] = 4'b1001;
	mem[1064] = 4'b1001;
	mem[1065] = 4'b1001;
	mem[1066] = 4'b1010;
	mem[1067] = 4'b1011;
	mem[1068] = 4'b1011;
	mem[1069] = 4'b1011;
	mem[1070] = 4'b1011;
	mem[1071] = 4'b1011;
	mem[1072] = 4'b1100;
	mem[1073] = 4'b1100;
	mem[1074] = 4'b1100;
	mem[1075] = 4'b1100;
	mem[1076] = 4'b1100;
	mem[1077] = 4'b1101;
	mem[1078] = 4'b1110;
	mem[1079] = 4'b1110;
	mem[1080] = 4'b1110;
	mem[1081] = 4'b1110;
	mem[1082] = 4'b1110;
	mem[1083] = 4'b1111;
	mem[1084] = 4'b1111;
	mem[1085] = 4'b1111;
	mem[1086] = 4'b1111;
	mem[1087] = 4'b1111;
	mem[1088] = 4'b1111;
	mem[1089] = 4'b1111;
	mem[1090] = 4'b1111;
	mem[1091] = 4'b1110;
	mem[1092] = 4'b1101;
	mem[1093] = 4'b1110;
	mem[1094] = 4'b0111;
	mem[1095] = 4'b0010;
	mem[1096] = 4'b0001;
	mem[1097] = 4'b0001;
	mem[1098] = 4'b0010;
	mem[1099] = 4'b0010;
	mem[1100] = 4'b0010;
	mem[1101] = 4'b0010;
	mem[1102] = 4'b0010;
	mem[1103] = 4'b0011;
	mem[1104] = 4'b0011;
	mem[1105] = 4'b0010;
	mem[1106] = 4'b0010;
	mem[1107] = 4'b0010;
	mem[1108] = 4'b0010;
	mem[1109] = 4'b0011;
	mem[1110] = 4'b0011;
	mem[1111] = 4'b0011;
	mem[1112] = 4'b0011;
	mem[1113] = 4'b0011;
	mem[1114] = 4'b0011;
	mem[1115] = 4'b0011;
	mem[1116] = 4'b0011;
	mem[1117] = 4'b0011;
	mem[1118] = 4'b0100;
	mem[1119] = 4'b0100;
	mem[1120] = 4'b0100;
	mem[1121] = 4'b0100;
	mem[1122] = 4'b0100;
	mem[1123] = 4'b0100;
	mem[1124] = 4'b0100;
	mem[1125] = 4'b0100;
	mem[1126] = 4'b0100;
	mem[1127] = 4'b0101;
	mem[1128] = 4'b0101;
	mem[1129] = 4'b0101;
	mem[1130] = 4'b0101;
	mem[1131] = 4'b0101;
	mem[1132] = 4'b0101;
	mem[1133] = 4'b0101;
	mem[1134] = 4'b0101;
	mem[1135] = 4'b0101;
	mem[1136] = 4'b0101;
	mem[1137] = 4'b0110;
	mem[1138] = 4'b0110;
	mem[1139] = 4'b0110;
	mem[1140] = 4'b0110;
	mem[1141] = 4'b0110;
	mem[1142] = 4'b0110;
	mem[1143] = 4'b0110;
	mem[1144] = 4'b0110;
	mem[1145] = 4'b0110;
	mem[1146] = 4'b0001;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0000;
	mem[1156] = 4'b0000;
	mem[1157] = 4'b0000;
	mem[1158] = 4'b0000;
	mem[1159] = 4'b0000;
	mem[1160] = 4'b0000;
	mem[1161] = 4'b0001;
	mem[1162] = 4'b0001;
	mem[1163] = 4'b0001;
	mem[1164] = 4'b0001;
	mem[1165] = 4'b0001;
	mem[1166] = 4'b0010;
	mem[1167] = 4'b0011;
	mem[1168] = 4'b0011;
	mem[1169] = 4'b0011;
	mem[1170] = 4'b0100;
	mem[1171] = 4'b0011;
	mem[1172] = 4'b0100;
	mem[1173] = 4'b0101;
	mem[1174] = 4'b0101;
	mem[1175] = 4'b0100;
	mem[1176] = 4'b0100;
	mem[1177] = 4'b0101;
	mem[1178] = 4'b0110;
	mem[1179] = 4'b0110;
	mem[1180] = 4'b0110;
	mem[1181] = 4'b0110;
	mem[1182] = 4'b0110;
	mem[1183] = 4'b0111;
	mem[1184] = 4'b1000;
	mem[1185] = 4'b1000;
	mem[1186] = 4'b1000;
	mem[1187] = 4'b1000;
	mem[1188] = 4'b1000;
	mem[1189] = 4'b1001;
	mem[1190] = 4'b1001;
	mem[1191] = 4'b1001;
	mem[1192] = 4'b1001;
	mem[1193] = 4'b1001;
	mem[1194] = 4'b1010;
	mem[1195] = 4'b1011;
	mem[1196] = 4'b1011;
	mem[1197] = 4'b1011;
	mem[1198] = 4'b1011;
	mem[1199] = 4'b1011;
	mem[1200] = 4'b1100;
	mem[1201] = 4'b1100;
	mem[1202] = 4'b1100;
	mem[1203] = 4'b1100;
	mem[1204] = 4'b1100;
	mem[1205] = 4'b1101;
	mem[1206] = 4'b1110;
	mem[1207] = 4'b1110;
	mem[1208] = 4'b1110;
	mem[1209] = 4'b1110;
	mem[1210] = 4'b1110;
	mem[1211] = 4'b1111;
	mem[1212] = 4'b1111;
	mem[1213] = 4'b1111;
	mem[1214] = 4'b1111;
	mem[1215] = 4'b1111;
	mem[1216] = 4'b1111;
	mem[1217] = 4'b1111;
	mem[1218] = 4'b1111;
	mem[1219] = 4'b1101;
	mem[1220] = 4'b1110;
	mem[1221] = 4'b1111;
	mem[1222] = 4'b0111;
	mem[1223] = 4'b0001;
	mem[1224] = 4'b0010;
	mem[1225] = 4'b0010;
	mem[1226] = 4'b0010;
	mem[1227] = 4'b0011;
	mem[1228] = 4'b0010;
	mem[1229] = 4'b0010;
	mem[1230] = 4'b0011;
	mem[1231] = 4'b0011;
	mem[1232] = 4'b0011;
	mem[1233] = 4'b0010;
	mem[1234] = 4'b0010;
	mem[1235] = 4'b0011;
	mem[1236] = 4'b0011;
	mem[1237] = 4'b0011;
	mem[1238] = 4'b0011;
	mem[1239] = 4'b0011;
	mem[1240] = 4'b0011;
	mem[1241] = 4'b0011;
	mem[1242] = 4'b0011;
	mem[1243] = 4'b0011;
	mem[1244] = 4'b0100;
	mem[1245] = 4'b0100;
	mem[1246] = 4'b0100;
	mem[1247] = 4'b0100;
	mem[1248] = 4'b0100;
	mem[1249] = 4'b0100;
	mem[1250] = 4'b0100;
	mem[1251] = 4'b0100;
	mem[1252] = 4'b0100;
	mem[1253] = 4'b0101;
	mem[1254] = 4'b0101;
	mem[1255] = 4'b0101;
	mem[1256] = 4'b0101;
	mem[1257] = 4'b0101;
	mem[1258] = 4'b0101;
	mem[1259] = 4'b0101;
	mem[1260] = 4'b0101;
	mem[1261] = 4'b0101;
	mem[1262] = 4'b0110;
	mem[1263] = 4'b0110;
	mem[1264] = 4'b0110;
	mem[1265] = 4'b0110;
	mem[1266] = 4'b0110;
	mem[1267] = 4'b0110;
	mem[1268] = 4'b0110;
	mem[1269] = 4'b0110;
	mem[1270] = 4'b0110;
	mem[1271] = 4'b0111;
	mem[1272] = 4'b0111;
	mem[1273] = 4'b0110;
	mem[1274] = 4'b0001;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0000;
	mem[1284] = 4'b0000;
	mem[1285] = 4'b0000;
	mem[1286] = 4'b0000;
	mem[1287] = 4'b0000;
	mem[1288] = 4'b0000;
	mem[1289] = 4'b0001;
	mem[1290] = 4'b0001;
	mem[1291] = 4'b0001;
	mem[1292] = 4'b0001;
	mem[1293] = 4'b0001;
	mem[1294] = 4'b0010;
	mem[1295] = 4'b0011;
	mem[1296] = 4'b0011;
	mem[1297] = 4'b0100;
	mem[1298] = 4'b0011;
	mem[1299] = 4'b0011;
	mem[1300] = 4'b0100;
	mem[1301] = 4'b0100;
	mem[1302] = 4'b0100;
	mem[1303] = 4'b0100;
	mem[1304] = 4'b0100;
	mem[1305] = 4'b0101;
	mem[1306] = 4'b0110;
	mem[1307] = 4'b0101;
	mem[1308] = 4'b0110;
	mem[1309] = 4'b0110;
	mem[1310] = 4'b0110;
	mem[1311] = 4'b0111;
	mem[1312] = 4'b1000;
	mem[1313] = 4'b1000;
	mem[1314] = 4'b1000;
	mem[1315] = 4'b1000;
	mem[1316] = 4'b1000;
	mem[1317] = 4'b1001;
	mem[1318] = 4'b1001;
	mem[1319] = 4'b1001;
	mem[1320] = 4'b1001;
	mem[1321] = 4'b1001;
	mem[1322] = 4'b1010;
	mem[1323] = 4'b1011;
	mem[1324] = 4'b1011;
	mem[1325] = 4'b1011;
	mem[1326] = 4'b1011;
	mem[1327] = 4'b1011;
	mem[1328] = 4'b1100;
	mem[1329] = 4'b1100;
	mem[1330] = 4'b1100;
	mem[1331] = 4'b1100;
	mem[1332] = 4'b1100;
	mem[1333] = 4'b1101;
	mem[1334] = 4'b1110;
	mem[1335] = 4'b1110;
	mem[1336] = 4'b1110;
	mem[1337] = 4'b1110;
	mem[1338] = 4'b1110;
	mem[1339] = 4'b1111;
	mem[1340] = 4'b1111;
	mem[1341] = 4'b1111;
	mem[1342] = 4'b1111;
	mem[1343] = 4'b1111;
	mem[1344] = 4'b1111;
	mem[1345] = 4'b1111;
	mem[1346] = 4'b1110;
	mem[1347] = 4'b1101;
	mem[1348] = 4'b1110;
	mem[1349] = 4'b1111;
	mem[1350] = 4'b0111;
	mem[1351] = 4'b0010;
	mem[1352] = 4'b0010;
	mem[1353] = 4'b0010;
	mem[1354] = 4'b0010;
	mem[1355] = 4'b0011;
	mem[1356] = 4'b0011;
	mem[1357] = 4'b0010;
	mem[1358] = 4'b0010;
	mem[1359] = 4'b0011;
	mem[1360] = 4'b0011;
	mem[1361] = 4'b0011;
	mem[1362] = 4'b0011;
	mem[1363] = 4'b0011;
	mem[1364] = 4'b0011;
	mem[1365] = 4'b0011;
	mem[1366] = 4'b0011;
	mem[1367] = 4'b0011;
	mem[1368] = 4'b0011;
	mem[1369] = 4'b0100;
	mem[1370] = 4'b0100;
	mem[1371] = 4'b0100;
	mem[1372] = 4'b0100;
	mem[1373] = 4'b0100;
	mem[1374] = 4'b0100;
	mem[1375] = 4'b0100;
	mem[1376] = 4'b0100;
	mem[1377] = 4'b0100;
	mem[1378] = 4'b0101;
	mem[1379] = 4'b0101;
	mem[1380] = 4'b0101;
	mem[1381] = 4'b0101;
	mem[1382] = 4'b0101;
	mem[1383] = 4'b0101;
	mem[1384] = 4'b0101;
	mem[1385] = 4'b0101;
	mem[1386] = 4'b0101;
	mem[1387] = 4'b0110;
	mem[1388] = 4'b0110;
	mem[1389] = 4'b0110;
	mem[1390] = 4'b0110;
	mem[1391] = 4'b0110;
	mem[1392] = 4'b0110;
	mem[1393] = 4'b0110;
	mem[1394] = 4'b0110;
	mem[1395] = 4'b0110;
	mem[1396] = 4'b0110;
	mem[1397] = 4'b0111;
	mem[1398] = 4'b0111;
	mem[1399] = 4'b0111;
	mem[1400] = 4'b0111;
	mem[1401] = 4'b0111;
	mem[1402] = 4'b0001;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0000;
	mem[1412] = 4'b0000;
	mem[1413] = 4'b0000;
	mem[1414] = 4'b0000;
	mem[1415] = 4'b0000;
	mem[1416] = 4'b0000;
	mem[1417] = 4'b0001;
	mem[1418] = 4'b0001;
	mem[1419] = 4'b0001;
	mem[1420] = 4'b0001;
	mem[1421] = 4'b0001;
	mem[1422] = 4'b0010;
	mem[1423] = 4'b0011;
	mem[1424] = 4'b0011;
	mem[1425] = 4'b0100;
	mem[1426] = 4'b0011;
	mem[1427] = 4'b0011;
	mem[1428] = 4'b0100;
	mem[1429] = 4'b0100;
	mem[1430] = 4'b0100;
	mem[1431] = 4'b0100;
	mem[1432] = 4'b0100;
	mem[1433] = 4'b0101;
	mem[1434] = 4'b0101;
	mem[1435] = 4'b0101;
	mem[1436] = 4'b0110;
	mem[1437] = 4'b0110;
	mem[1438] = 4'b0110;
	mem[1439] = 4'b0111;
	mem[1440] = 4'b1000;
	mem[1441] = 4'b1000;
	mem[1442] = 4'b1000;
	mem[1443] = 4'b1000;
	mem[1444] = 4'b1000;
	mem[1445] = 4'b1001;
	mem[1446] = 4'b1001;
	mem[1447] = 4'b1001;
	mem[1448] = 4'b1001;
	mem[1449] = 4'b1001;
	mem[1450] = 4'b1010;
	mem[1451] = 4'b1011;
	mem[1452] = 4'b1011;
	mem[1453] = 4'b1011;
	mem[1454] = 4'b1011;
	mem[1455] = 4'b1011;
	mem[1456] = 4'b1100;
	mem[1457] = 4'b1100;
	mem[1458] = 4'b1100;
	mem[1459] = 4'b1100;
	mem[1460] = 4'b1100;
	mem[1461] = 4'b1101;
	mem[1462] = 4'b1110;
	mem[1463] = 4'b1110;
	mem[1464] = 4'b1110;
	mem[1465] = 4'b1110;
	mem[1466] = 4'b1110;
	mem[1467] = 4'b1111;
	mem[1468] = 4'b1111;
	mem[1469] = 4'b1111;
	mem[1470] = 4'b1111;
	mem[1471] = 4'b1111;
	mem[1472] = 4'b1111;
	mem[1473] = 4'b1111;
	mem[1474] = 4'b1110;
	mem[1475] = 4'b1101;
	mem[1476] = 4'b1110;
	mem[1477] = 4'b1111;
	mem[1478] = 4'b0111;
	mem[1479] = 4'b0010;
	mem[1480] = 4'b0010;
	mem[1481] = 4'b0010;
	mem[1482] = 4'b0010;
	mem[1483] = 4'b0011;
	mem[1484] = 4'b0011;
	mem[1485] = 4'b0011;
	mem[1486] = 4'b0011;
	mem[1487] = 4'b0011;
	mem[1488] = 4'b0011;
	mem[1489] = 4'b0011;
	mem[1490] = 4'b0011;
	mem[1491] = 4'b0011;
	mem[1492] = 4'b0011;
	mem[1493] = 4'b0011;
	mem[1494] = 4'b0011;
	mem[1495] = 4'b0100;
	mem[1496] = 4'b0100;
	mem[1497] = 4'b0100;
	mem[1498] = 4'b0100;
	mem[1499] = 4'b0100;
	mem[1500] = 4'b0100;
	mem[1501] = 4'b0100;
	mem[1502] = 4'b0100;
	mem[1503] = 4'b0100;
	mem[1504] = 4'b0101;
	mem[1505] = 4'b0101;
	mem[1506] = 4'b0101;
	mem[1507] = 4'b0101;
	mem[1508] = 4'b0101;
	mem[1509] = 4'b0101;
	mem[1510] = 4'b0101;
	mem[1511] = 4'b0101;
	mem[1512] = 4'b0101;
	mem[1513] = 4'b0110;
	mem[1514] = 4'b0110;
	mem[1515] = 4'b0110;
	mem[1516] = 4'b0110;
	mem[1517] = 4'b0110;
	mem[1518] = 4'b0110;
	mem[1519] = 4'b0110;
	mem[1520] = 4'b0110;
	mem[1521] = 4'b0110;
	mem[1522] = 4'b0111;
	mem[1523] = 4'b0111;
	mem[1524] = 4'b0111;
	mem[1525] = 4'b0111;
	mem[1526] = 4'b0111;
	mem[1527] = 4'b0111;
	mem[1528] = 4'b0111;
	mem[1529] = 4'b0111;
	mem[1530] = 4'b0001;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0000;
	mem[1540] = 4'b0000;
	mem[1541] = 4'b0000;
	mem[1542] = 4'b0000;
	mem[1543] = 4'b0000;
	mem[1544] = 4'b0000;
	mem[1545] = 4'b0001;
	mem[1546] = 4'b0001;
	mem[1547] = 4'b0001;
	mem[1548] = 4'b0001;
	mem[1549] = 4'b0001;
	mem[1550] = 4'b0010;
	mem[1551] = 4'b0010;
	mem[1552] = 4'b0010;
	mem[1553] = 4'b0011;
	mem[1554] = 4'b0010;
	mem[1555] = 4'b0010;
	mem[1556] = 4'b0100;
	mem[1557] = 4'b0100;
	mem[1558] = 4'b0100;
	mem[1559] = 4'b0100;
	mem[1560] = 4'b0100;
	mem[1561] = 4'b0100;
	mem[1562] = 4'b0101;
	mem[1563] = 4'b0101;
	mem[1564] = 4'b0101;
	mem[1565] = 4'b0110;
	mem[1566] = 4'b0101;
	mem[1567] = 4'b0110;
	mem[1568] = 4'b0111;
	mem[1569] = 4'b0111;
	mem[1570] = 4'b0111;
	mem[1571] = 4'b0111;
	mem[1572] = 4'b0111;
	mem[1573] = 4'b1000;
	mem[1574] = 4'b1000;
	mem[1575] = 4'b1000;
	mem[1576] = 4'b1000;
	mem[1577] = 4'b1000;
	mem[1578] = 4'b1001;
	mem[1579] = 4'b1010;
	mem[1580] = 4'b1010;
	mem[1581] = 4'b1010;
	mem[1582] = 4'b1010;
	mem[1583] = 4'b1010;
	mem[1584] = 4'b1011;
	mem[1585] = 4'b1011;
	mem[1586] = 4'b1011;
	mem[1587] = 4'b1011;
	mem[1588] = 4'b1011;
	mem[1589] = 4'b1100;
	mem[1590] = 4'b1101;
	mem[1591] = 4'b1101;
	mem[1592] = 4'b1101;
	mem[1593] = 4'b1101;
	mem[1594] = 4'b1101;
	mem[1595] = 4'b1101;
	mem[1596] = 4'b1101;
	mem[1597] = 4'b1101;
	mem[1598] = 4'b1101;
	mem[1599] = 4'b1101;
	mem[1600] = 4'b1101;
	mem[1601] = 4'b1110;
	mem[1602] = 4'b1110;
	mem[1603] = 4'b1100;
	mem[1604] = 4'b1100;
	mem[1605] = 4'b1101;
	mem[1606] = 4'b0111;
	mem[1607] = 4'b0010;
	mem[1608] = 4'b0010;
	mem[1609] = 4'b0010;
	mem[1610] = 4'b0010;
	mem[1611] = 4'b0011;
	mem[1612] = 4'b0011;
	mem[1613] = 4'b0010;
	mem[1614] = 4'b0011;
	mem[1615] = 4'b0011;
	mem[1616] = 4'b0011;
	mem[1617] = 4'b0011;
	mem[1618] = 4'b0011;
	mem[1619] = 4'b0011;
	mem[1620] = 4'b0011;
	mem[1621] = 4'b0011;
	mem[1622] = 4'b0011;
	mem[1623] = 4'b0011;
	mem[1624] = 4'b0100;
	mem[1625] = 4'b0100;
	mem[1626] = 4'b0100;
	mem[1627] = 4'b0100;
	mem[1628] = 4'b0100;
	mem[1629] = 4'b0100;
	mem[1630] = 4'b0100;
	mem[1631] = 4'b0100;
	mem[1632] = 4'b0100;
	mem[1633] = 4'b0100;
	mem[1634] = 4'b0101;
	mem[1635] = 4'b0101;
	mem[1636] = 4'b0101;
	mem[1637] = 4'b0101;
	mem[1638] = 4'b0101;
	mem[1639] = 4'b0101;
	mem[1640] = 4'b0101;
	mem[1641] = 4'b0101;
	mem[1642] = 4'b0101;
	mem[1643] = 4'b0101;
	mem[1644] = 4'b0110;
	mem[1645] = 4'b0110;
	mem[1646] = 4'b0110;
	mem[1647] = 4'b0110;
	mem[1648] = 4'b0110;
	mem[1649] = 4'b0110;
	mem[1650] = 4'b0110;
	mem[1651] = 4'b0110;
	mem[1652] = 4'b0110;
	mem[1653] = 4'b0110;
	mem[1654] = 4'b0111;
	mem[1655] = 4'b0111;
	mem[1656] = 4'b0111;
	mem[1657] = 4'b0111;
	mem[1658] = 4'b0001;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0000;
	mem[1668] = 4'b0000;
	mem[1669] = 4'b0000;
	mem[1670] = 4'b0000;
	mem[1671] = 4'b0000;
	mem[1672] = 4'b0000;
	mem[1673] = 4'b0000;
	mem[1674] = 4'b0000;
	mem[1675] = 4'b0000;
	mem[1676] = 4'b0000;
	mem[1677] = 4'b0000;
	mem[1678] = 4'b0000;
	mem[1679] = 4'b0000;
	mem[1680] = 4'b0000;
	mem[1681] = 4'b0001;
	mem[1682] = 4'b0000;
	mem[1683] = 4'b0000;
	mem[1684] = 4'b0000;
	mem[1685] = 4'b0000;
	mem[1686] = 4'b0000;
	mem[1687] = 4'b0000;
	mem[1688] = 4'b0000;
	mem[1689] = 4'b0001;
	mem[1690] = 4'b0000;
	mem[1691] = 4'b0001;
	mem[1692] = 4'b0001;
	mem[1693] = 4'b0001;
	mem[1694] = 4'b0000;
	mem[1695] = 4'b0000;
	mem[1696] = 4'b0000;
	mem[1697] = 4'b0000;
	mem[1698] = 4'b0000;
	mem[1699] = 4'b0000;
	mem[1700] = 4'b0000;
	mem[1701] = 4'b0000;
	mem[1702] = 4'b0000;
	mem[1703] = 4'b0000;
	mem[1704] = 4'b0000;
	mem[1705] = 4'b0000;
	mem[1706] = 4'b0000;
	mem[1707] = 4'b0001;
	mem[1708] = 4'b0001;
	mem[1709] = 4'b0001;
	mem[1710] = 4'b0001;
	mem[1711] = 4'b0001;
	mem[1712] = 4'b0001;
	mem[1713] = 4'b0001;
	mem[1714] = 4'b0001;
	mem[1715] = 4'b0001;
	mem[1716] = 4'b0001;
	mem[1717] = 4'b0001;
	mem[1718] = 4'b0001;
	mem[1719] = 4'b0001;
	mem[1720] = 4'b0001;
	mem[1721] = 4'b0001;
	mem[1722] = 4'b0001;
	mem[1723] = 4'b0001;
	mem[1724] = 4'b0001;
	mem[1725] = 4'b0001;
	mem[1726] = 4'b0001;
	mem[1727] = 4'b0001;
	mem[1728] = 4'b0001;
	mem[1729] = 4'b0010;
	mem[1730] = 4'b0001;
	mem[1731] = 4'b0010;
	mem[1732] = 4'b0001;
	mem[1733] = 4'b0001;
	mem[1734] = 4'b0001;
	mem[1735] = 4'b0000;
	mem[1736] = 4'b0000;
	mem[1737] = 4'b0000;
	mem[1738] = 4'b0001;
	mem[1739] = 4'b0001;
	mem[1740] = 4'b0000;
	mem[1741] = 4'b0000;
	mem[1742] = 4'b0000;
	mem[1743] = 4'b0000;
	mem[1744] = 4'b0000;
	mem[1745] = 4'b0000;
	mem[1746] = 4'b0000;
	mem[1747] = 4'b0000;
	mem[1748] = 4'b0000;
	mem[1749] = 4'b0000;
	mem[1750] = 4'b0000;
	mem[1751] = 4'b0000;
	mem[1752] = 4'b0000;
	mem[1753] = 4'b0000;
	mem[1754] = 4'b0000;
	mem[1755] = 4'b0000;
	mem[1756] = 4'b0000;
	mem[1757] = 4'b0000;
	mem[1758] = 4'b0000;
	mem[1759] = 4'b0000;
	mem[1760] = 4'b0000;
	mem[1761] = 4'b0000;
	mem[1762] = 4'b0000;
	mem[1763] = 4'b0000;
	mem[1764] = 4'b0000;
	mem[1765] = 4'b0000;
	mem[1766] = 4'b0000;
	mem[1767] = 4'b0000;
	mem[1768] = 4'b0000;
	mem[1769] = 4'b0000;
	mem[1770] = 4'b0000;
	mem[1771] = 4'b0000;
	mem[1772] = 4'b0000;
	mem[1773] = 4'b0000;
	mem[1774] = 4'b0000;
	mem[1775] = 4'b0000;
	mem[1776] = 4'b0000;
	mem[1777] = 4'b0000;
	mem[1778] = 4'b0000;
	mem[1779] = 4'b0000;
	mem[1780] = 4'b0000;
	mem[1781] = 4'b0000;
	mem[1782] = 4'b0000;
	mem[1783] = 4'b0000;
	mem[1784] = 4'b0000;
	mem[1785] = 4'b0000;
	mem[1786] = 4'b0000;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0000;
	mem[1796] = 4'b0000;
	mem[1797] = 4'b0000;
	mem[1798] = 4'b0000;
	mem[1799] = 4'b0000;
	mem[1800] = 4'b0000;
	mem[1801] = 4'b0000;
	mem[1802] = 4'b0000;
	mem[1803] = 4'b0000;
	mem[1804] = 4'b0000;
	mem[1805] = 4'b0000;
	mem[1806] = 4'b0000;
	mem[1807] = 4'b0000;
	mem[1808] = 4'b0000;
	mem[1809] = 4'b0000;
	mem[1810] = 4'b0001;
	mem[1811] = 4'b0000;
	mem[1812] = 4'b0000;
	mem[1813] = 4'b0000;
	mem[1814] = 4'b0000;
	mem[1815] = 4'b0000;
	mem[1816] = 4'b0000;
	mem[1817] = 4'b0000;
	mem[1818] = 4'b0000;
	mem[1819] = 4'b0000;
	mem[1820] = 4'b0000;
	mem[1821] = 4'b0001;
	mem[1822] = 4'b0000;
	mem[1823] = 4'b0000;
	mem[1824] = 4'b0000;
	mem[1825] = 4'b0000;
	mem[1826] = 4'b0000;
	mem[1827] = 4'b0000;
	mem[1828] = 4'b0000;
	mem[1829] = 4'b0000;
	mem[1830] = 4'b0000;
	mem[1831] = 4'b0000;
	mem[1832] = 4'b0000;
	mem[1833] = 4'b0000;
	mem[1834] = 4'b0000;
	mem[1835] = 4'b0000;
	mem[1836] = 4'b0000;
	mem[1837] = 4'b0000;
	mem[1838] = 4'b0000;
	mem[1839] = 4'b0000;
	mem[1840] = 4'b0000;
	mem[1841] = 4'b0000;
	mem[1842] = 4'b0000;
	mem[1843] = 4'b0000;
	mem[1844] = 4'b0000;
	mem[1845] = 4'b0000;
	mem[1846] = 4'b0000;
	mem[1847] = 4'b0000;
	mem[1848] = 4'b0000;
	mem[1849] = 4'b0000;
	mem[1850] = 4'b0000;
	mem[1851] = 4'b0000;
	mem[1852] = 4'b0000;
	mem[1853] = 4'b0000;
	mem[1854] = 4'b0000;
	mem[1855] = 4'b0000;
	mem[1856] = 4'b0000;
	mem[1857] = 4'b0001;
	mem[1858] = 4'b0000;
	mem[1859] = 4'b0000;
	mem[1860] = 4'b0000;
	mem[1861] = 4'b0000;
	mem[1862] = 4'b0000;
	mem[1863] = 4'b0000;
	mem[1864] = 4'b0000;
	mem[1865] = 4'b0001;
	mem[1866] = 4'b0001;
	mem[1867] = 4'b0000;
	mem[1868] = 4'b0000;
	mem[1869] = 4'b0000;
	mem[1870] = 4'b0000;
	mem[1871] = 4'b0000;
	mem[1872] = 4'b0000;
	mem[1873] = 4'b0000;
	mem[1874] = 4'b0000;
	mem[1875] = 4'b0000;
	mem[1876] = 4'b0000;
	mem[1877] = 4'b0000;
	mem[1878] = 4'b0000;
	mem[1879] = 4'b0000;
	mem[1880] = 4'b0000;
	mem[1881] = 4'b0000;
	mem[1882] = 4'b0000;
	mem[1883] = 4'b0000;
	mem[1884] = 4'b0000;
	mem[1885] = 4'b0000;
	mem[1886] = 4'b0000;
	mem[1887] = 4'b0000;
	mem[1888] = 4'b0000;
	mem[1889] = 4'b0000;
	mem[1890] = 4'b0000;
	mem[1891] = 4'b0000;
	mem[1892] = 4'b0000;
	mem[1893] = 4'b0000;
	mem[1894] = 4'b0000;
	mem[1895] = 4'b0000;
	mem[1896] = 4'b0000;
	mem[1897] = 4'b0000;
	mem[1898] = 4'b0000;
	mem[1899] = 4'b0000;
	mem[1900] = 4'b0000;
	mem[1901] = 4'b0000;
	mem[1902] = 4'b0000;
	mem[1903] = 4'b0000;
	mem[1904] = 4'b0000;
	mem[1905] = 4'b0000;
	mem[1906] = 4'b0000;
	mem[1907] = 4'b0000;
	mem[1908] = 4'b0000;
	mem[1909] = 4'b0000;
	mem[1910] = 4'b0000;
	mem[1911] = 4'b0000;
	mem[1912] = 4'b0000;
	mem[1913] = 4'b0000;
	mem[1914] = 4'b0000;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0000;
	mem[1924] = 4'b0000;
	mem[1925] = 4'b0000;
	mem[1926] = 4'b0000;
	mem[1927] = 4'b0000;
	mem[1928] = 4'b0000;
	mem[1929] = 4'b0000;
	mem[1930] = 4'b0000;
	mem[1931] = 4'b0000;
	mem[1932] = 4'b0000;
	mem[1933] = 4'b0000;
	mem[1934] = 4'b0000;
	mem[1935] = 4'b0000;
	mem[1936] = 4'b0000;
	mem[1937] = 4'b0000;
	mem[1938] = 4'b0000;
	mem[1939] = 4'b0000;
	mem[1940] = 4'b0000;
	mem[1941] = 4'b0000;
	mem[1942] = 4'b0000;
	mem[1943] = 4'b0000;
	mem[1944] = 4'b0000;
	mem[1945] = 4'b0000;
	mem[1946] = 4'b0000;
	mem[1947] = 4'b0000;
	mem[1948] = 4'b0001;
	mem[1949] = 4'b0000;
	mem[1950] = 4'b0000;
	mem[1951] = 4'b0000;
	mem[1952] = 4'b0000;
	mem[1953] = 4'b0000;
	mem[1954] = 4'b0000;
	mem[1955] = 4'b0000;
	mem[1956] = 4'b0000;
	mem[1957] = 4'b0000;
	mem[1958] = 4'b0000;
	mem[1959] = 4'b0000;
	mem[1960] = 4'b0000;
	mem[1961] = 4'b0000;
	mem[1962] = 4'b0000;
	mem[1963] = 4'b0000;
	mem[1964] = 4'b0000;
	mem[1965] = 4'b0000;
	mem[1966] = 4'b0000;
	mem[1967] = 4'b0000;
	mem[1968] = 4'b0000;
	mem[1969] = 4'b0000;
	mem[1970] = 4'b0000;
	mem[1971] = 4'b0000;
	mem[1972] = 4'b0000;
	mem[1973] = 4'b0000;
	mem[1974] = 4'b0000;
	mem[1975] = 4'b0000;
	mem[1976] = 4'b0000;
	mem[1977] = 4'b0000;
	mem[1978] = 4'b0000;
	mem[1979] = 4'b0000;
	mem[1980] = 4'b0000;
	mem[1981] = 4'b0000;
	mem[1982] = 4'b0001;
	mem[1983] = 4'b0001;
	mem[1984] = 4'b0001;
	mem[1985] = 4'b0000;
	mem[1986] = 4'b0000;
	mem[1987] = 4'b0000;
	mem[1988] = 4'b0000;
	mem[1989] = 4'b0000;
	mem[1990] = 4'b0001;
	mem[1991] = 4'b0001;
	mem[1992] = 4'b0001;
	mem[1993] = 4'b0001;
	mem[1994] = 4'b0000;
	mem[1995] = 4'b0000;
	mem[1996] = 4'b0000;
	mem[1997] = 4'b0000;
	mem[1998] = 4'b0000;
	mem[1999] = 4'b0000;
	mem[2000] = 4'b0000;
	mem[2001] = 4'b0000;
	mem[2002] = 4'b0000;
	mem[2003] = 4'b0000;
	mem[2004] = 4'b0000;
	mem[2005] = 4'b0000;
	mem[2006] = 4'b0000;
	mem[2007] = 4'b0000;
	mem[2008] = 4'b0000;
	mem[2009] = 4'b0000;
	mem[2010] = 4'b0000;
	mem[2011] = 4'b0000;
	mem[2012] = 4'b0000;
	mem[2013] = 4'b0000;
	mem[2014] = 4'b0000;
	mem[2015] = 4'b0000;
	mem[2016] = 4'b0000;
	mem[2017] = 4'b0000;
	mem[2018] = 4'b0000;
	mem[2019] = 4'b0000;
	mem[2020] = 4'b0000;
	mem[2021] = 4'b0000;
	mem[2022] = 4'b0000;
	mem[2023] = 4'b0000;
	mem[2024] = 4'b0000;
	mem[2025] = 4'b0000;
	mem[2026] = 4'b0000;
	mem[2027] = 4'b0000;
	mem[2028] = 4'b0000;
	mem[2029] = 4'b0000;
	mem[2030] = 4'b0000;
	mem[2031] = 4'b0000;
	mem[2032] = 4'b0000;
	mem[2033] = 4'b0000;
	mem[2034] = 4'b0000;
	mem[2035] = 4'b0000;
	mem[2036] = 4'b0000;
	mem[2037] = 4'b0000;
	mem[2038] = 4'b0000;
	mem[2039] = 4'b0000;
	mem[2040] = 4'b0000;
	mem[2041] = 4'b0000;
	mem[2042] = 4'b0000;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0000;
	mem[2052] = 4'b0000;
	mem[2053] = 4'b0000;
	mem[2054] = 4'b0000;
	mem[2055] = 4'b0000;
	mem[2056] = 4'b0000;
	mem[2057] = 4'b0000;
	mem[2058] = 4'b0000;
	mem[2059] = 4'b0000;
	mem[2060] = 4'b0000;
	mem[2061] = 4'b0000;
	mem[2062] = 4'b0000;
	mem[2063] = 4'b0000;
	mem[2064] = 4'b0000;
	mem[2065] = 4'b0000;
	mem[2066] = 4'b0000;
	mem[2067] = 4'b0000;
	mem[2068] = 4'b0000;
	mem[2069] = 4'b0000;
	mem[2070] = 4'b0000;
	mem[2071] = 4'b0000;
	mem[2072] = 4'b0000;
	mem[2073] = 4'b0000;
	mem[2074] = 4'b0000;
	mem[2075] = 4'b0000;
	mem[2076] = 4'b0001;
	mem[2077] = 4'b0000;
	mem[2078] = 4'b0000;
	mem[2079] = 4'b0000;
	mem[2080] = 4'b0000;
	mem[2081] = 4'b0000;
	mem[2082] = 4'b0000;
	mem[2083] = 4'b0000;
	mem[2084] = 4'b0000;
	mem[2085] = 4'b0000;
	mem[2086] = 4'b0000;
	mem[2087] = 4'b0000;
	mem[2088] = 4'b0000;
	mem[2089] = 4'b0000;
	mem[2090] = 4'b0000;
	mem[2091] = 4'b0000;
	mem[2092] = 4'b0000;
	mem[2093] = 4'b0000;
	mem[2094] = 4'b0000;
	mem[2095] = 4'b0000;
	mem[2096] = 4'b0000;
	mem[2097] = 4'b0000;
	mem[2098] = 4'b0000;
	mem[2099] = 4'b0000;
	mem[2100] = 4'b0000;
	mem[2101] = 4'b0000;
	mem[2102] = 4'b0000;
	mem[2103] = 4'b0000;
	mem[2104] = 4'b0000;
	mem[2105] = 4'b0000;
	mem[2106] = 4'b0000;
	mem[2107] = 4'b0000;
	mem[2108] = 4'b0000;
	mem[2109] = 4'b0000;
	mem[2110] = 4'b0001;
	mem[2111] = 4'b0000;
	mem[2112] = 4'b0000;
	mem[2113] = 4'b0000;
	mem[2114] = 4'b0000;
	mem[2115] = 4'b0000;
	mem[2116] = 4'b0000;
	mem[2117] = 4'b0000;
	mem[2118] = 4'b0000;
	mem[2119] = 4'b0000;
	mem[2120] = 4'b0000;
	mem[2121] = 4'b0000;
	mem[2122] = 4'b0000;
	mem[2123] = 4'b0000;
	mem[2124] = 4'b0000;
	mem[2125] = 4'b0000;
	mem[2126] = 4'b0000;
	mem[2127] = 4'b0000;
	mem[2128] = 4'b0000;
	mem[2129] = 4'b0000;
	mem[2130] = 4'b0000;
	mem[2131] = 4'b0000;
	mem[2132] = 4'b0000;
	mem[2133] = 4'b0000;
	mem[2134] = 4'b0000;
	mem[2135] = 4'b0000;
	mem[2136] = 4'b0000;
	mem[2137] = 4'b0000;
	mem[2138] = 4'b0000;
	mem[2139] = 4'b0000;
	mem[2140] = 4'b0000;
	mem[2141] = 4'b0000;
	mem[2142] = 4'b0000;
	mem[2143] = 4'b0000;
	mem[2144] = 4'b0000;
	mem[2145] = 4'b0000;
	mem[2146] = 4'b0000;
	mem[2147] = 4'b0000;
	mem[2148] = 4'b0000;
	mem[2149] = 4'b0000;
	mem[2150] = 4'b0000;
	mem[2151] = 4'b0000;
	mem[2152] = 4'b0000;
	mem[2153] = 4'b0000;
	mem[2154] = 4'b0000;
	mem[2155] = 4'b0000;
	mem[2156] = 4'b0000;
	mem[2157] = 4'b0000;
	mem[2158] = 4'b0000;
	mem[2159] = 4'b0000;
	mem[2160] = 4'b0000;
	mem[2161] = 4'b0000;
	mem[2162] = 4'b0000;
	mem[2163] = 4'b0000;
	mem[2164] = 4'b0000;
	mem[2165] = 4'b0000;
	mem[2166] = 4'b0000;
	mem[2167] = 4'b0000;
	mem[2168] = 4'b0000;
	mem[2169] = 4'b0000;
	mem[2170] = 4'b0000;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0000;
	mem[2180] = 4'b0000;
	mem[2181] = 4'b0000;
	mem[2182] = 4'b0000;
	mem[2183] = 4'b0000;
	mem[2184] = 4'b0000;
	mem[2185] = 4'b0000;
	mem[2186] = 4'b0000;
	mem[2187] = 4'b0000;
	mem[2188] = 4'b0000;
	mem[2189] = 4'b0000;
	mem[2190] = 4'b0000;
	mem[2191] = 4'b0000;
	mem[2192] = 4'b0000;
	mem[2193] = 4'b0000;
	mem[2194] = 4'b0000;
	mem[2195] = 4'b0000;
	mem[2196] = 4'b0000;
	mem[2197] = 4'b0000;
	mem[2198] = 4'b0000;
	mem[2199] = 4'b0000;
	mem[2200] = 4'b0000;
	mem[2201] = 4'b0000;
	mem[2202] = 4'b0000;
	mem[2203] = 4'b0001;
	mem[2204] = 4'b0000;
	mem[2205] = 4'b0000;
	mem[2206] = 4'b0000;
	mem[2207] = 4'b0000;
	mem[2208] = 4'b0000;
	mem[2209] = 4'b0000;
	mem[2210] = 4'b0000;
	mem[2211] = 4'b0000;
	mem[2212] = 4'b0000;
	mem[2213] = 4'b0000;
	mem[2214] = 4'b0000;
	mem[2215] = 4'b0000;
	mem[2216] = 4'b0000;
	mem[2217] = 4'b0000;
	mem[2218] = 4'b0000;
	mem[2219] = 4'b0000;
	mem[2220] = 4'b0000;
	mem[2221] = 4'b0000;
	mem[2222] = 4'b0000;
	mem[2223] = 4'b0000;
	mem[2224] = 4'b0000;
	mem[2225] = 4'b0000;
	mem[2226] = 4'b0000;
	mem[2227] = 4'b0000;
	mem[2228] = 4'b0000;
	mem[2229] = 4'b0000;
	mem[2230] = 4'b0000;
	mem[2231] = 4'b0000;
	mem[2232] = 4'b0000;
	mem[2233] = 4'b0000;
	mem[2234] = 4'b0000;
	mem[2235] = 4'b0000;
	mem[2236] = 4'b0000;
	mem[2237] = 4'b0000;
	mem[2238] = 4'b0001;
	mem[2239] = 4'b0000;
	mem[2240] = 4'b0000;
	mem[2241] = 4'b0000;
	mem[2242] = 4'b0000;
	mem[2243] = 4'b0000;
	mem[2244] = 4'b0000;
	mem[2245] = 4'b0000;
	mem[2246] = 4'b0000;
	mem[2247] = 4'b0000;
	mem[2248] = 4'b0000;
	mem[2249] = 4'b0000;
	mem[2250] = 4'b0000;
	mem[2251] = 4'b0000;
	mem[2252] = 4'b0000;
	mem[2253] = 4'b0000;
	mem[2254] = 4'b0000;
	mem[2255] = 4'b0000;
	mem[2256] = 4'b0000;
	mem[2257] = 4'b0000;
	mem[2258] = 4'b0000;
	mem[2259] = 4'b0000;
	mem[2260] = 4'b0000;
	mem[2261] = 4'b0000;
	mem[2262] = 4'b0000;
	mem[2263] = 4'b0000;
	mem[2264] = 4'b0000;
	mem[2265] = 4'b0000;
	mem[2266] = 4'b0000;
	mem[2267] = 4'b0000;
	mem[2268] = 4'b0000;
	mem[2269] = 4'b0000;
	mem[2270] = 4'b0000;
	mem[2271] = 4'b0000;
	mem[2272] = 4'b0000;
	mem[2273] = 4'b0000;
	mem[2274] = 4'b0000;
	mem[2275] = 4'b0000;
	mem[2276] = 4'b0000;
	mem[2277] = 4'b0000;
	mem[2278] = 4'b0000;
	mem[2279] = 4'b0000;
	mem[2280] = 4'b0000;
	mem[2281] = 4'b0000;
	mem[2282] = 4'b0000;
	mem[2283] = 4'b0000;
	mem[2284] = 4'b0000;
	mem[2285] = 4'b0000;
	mem[2286] = 4'b0000;
	mem[2287] = 4'b0000;
	mem[2288] = 4'b0000;
	mem[2289] = 4'b0000;
	mem[2290] = 4'b0000;
	mem[2291] = 4'b0000;
	mem[2292] = 4'b0000;
	mem[2293] = 4'b0000;
	mem[2294] = 4'b0000;
	mem[2295] = 4'b0000;
	mem[2296] = 4'b0000;
	mem[2297] = 4'b0000;
	mem[2298] = 4'b0000;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0000;
	mem[2308] = 4'b0000;
	mem[2309] = 4'b0000;
	mem[2310] = 4'b0000;
	mem[2311] = 4'b0000;
	mem[2312] = 4'b0000;
	mem[2313] = 4'b0000;
	mem[2314] = 4'b0000;
	mem[2315] = 4'b0000;
	mem[2316] = 4'b0000;
	mem[2317] = 4'b0000;
	mem[2318] = 4'b0000;
	mem[2319] = 4'b0000;
	mem[2320] = 4'b0000;
	mem[2321] = 4'b0000;
	mem[2322] = 4'b0000;
	mem[2323] = 4'b0000;
	mem[2324] = 4'b0000;
	mem[2325] = 4'b0000;
	mem[2326] = 4'b0000;
	mem[2327] = 4'b0000;
	mem[2328] = 4'b0000;
	mem[2329] = 4'b0000;
	mem[2330] = 4'b0001;
	mem[2331] = 4'b0001;
	mem[2332] = 4'b0000;
	mem[2333] = 4'b0000;
	mem[2334] = 4'b0000;
	mem[2335] = 4'b0000;
	mem[2336] = 4'b0000;
	mem[2337] = 4'b0000;
	mem[2338] = 4'b0000;
	mem[2339] = 4'b0000;
	mem[2340] = 4'b0000;
	mem[2341] = 4'b0000;
	mem[2342] = 4'b0000;
	mem[2343] = 4'b0000;
	mem[2344] = 4'b0000;
	mem[2345] = 4'b0000;
	mem[2346] = 4'b0000;
	mem[2347] = 4'b0000;
	mem[2348] = 4'b0000;
	mem[2349] = 4'b0000;
	mem[2350] = 4'b0000;
	mem[2351] = 4'b0000;
	mem[2352] = 4'b0000;
	mem[2353] = 4'b0000;
	mem[2354] = 4'b0000;
	mem[2355] = 4'b0000;
	mem[2356] = 4'b0000;
	mem[2357] = 4'b0000;
	mem[2358] = 4'b0000;
	mem[2359] = 4'b0000;
	mem[2360] = 4'b0000;
	mem[2361] = 4'b0000;
	mem[2362] = 4'b0000;
	mem[2363] = 4'b0000;
	mem[2364] = 4'b0000;
	mem[2365] = 4'b0000;
	mem[2366] = 4'b0000;
	mem[2367] = 4'b0000;
	mem[2368] = 4'b0000;
	mem[2369] = 4'b0000;
	mem[2370] = 4'b0000;
	mem[2371] = 4'b0000;
	mem[2372] = 4'b0001;
	mem[2373] = 4'b0000;
	mem[2374] = 4'b0000;
	mem[2375] = 4'b0000;
	mem[2376] = 4'b0000;
	mem[2377] = 4'b0000;
	mem[2378] = 4'b0000;
	mem[2379] = 4'b0000;
	mem[2380] = 4'b0000;
	mem[2381] = 4'b0000;
	mem[2382] = 4'b0000;
	mem[2383] = 4'b0000;
	mem[2384] = 4'b0000;
	mem[2385] = 4'b0000;
	mem[2386] = 4'b0000;
	mem[2387] = 4'b0000;
	mem[2388] = 4'b0000;
	mem[2389] = 4'b0000;
	mem[2390] = 4'b0000;
	mem[2391] = 4'b0000;
	mem[2392] = 4'b0000;
	mem[2393] = 4'b0000;
	mem[2394] = 4'b0000;
	mem[2395] = 4'b0000;
	mem[2396] = 4'b0000;
	mem[2397] = 4'b0000;
	mem[2398] = 4'b0000;
	mem[2399] = 4'b0000;
	mem[2400] = 4'b0000;
	mem[2401] = 4'b0000;
	mem[2402] = 4'b0000;
	mem[2403] = 4'b0000;
	mem[2404] = 4'b0000;
	mem[2405] = 4'b0000;
	mem[2406] = 4'b0000;
	mem[2407] = 4'b0000;
	mem[2408] = 4'b0000;
	mem[2409] = 4'b0000;
	mem[2410] = 4'b0000;
	mem[2411] = 4'b0000;
	mem[2412] = 4'b0000;
	mem[2413] = 4'b0000;
	mem[2414] = 4'b0000;
	mem[2415] = 4'b0000;
	mem[2416] = 4'b0000;
	mem[2417] = 4'b0000;
	mem[2418] = 4'b0000;
	mem[2419] = 4'b0000;
	mem[2420] = 4'b0000;
	mem[2421] = 4'b0000;
	mem[2422] = 4'b0000;
	mem[2423] = 4'b0000;
	mem[2424] = 4'b0000;
	mem[2425] = 4'b0000;
	mem[2426] = 4'b0000;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0000;
	mem[2436] = 4'b0000;
	mem[2437] = 4'b0000;
	mem[2438] = 4'b0000;
	mem[2439] = 4'b0000;
	mem[2440] = 4'b0000;
	mem[2441] = 4'b0000;
	mem[2442] = 4'b0000;
	mem[2443] = 4'b0000;
	mem[2444] = 4'b0000;
	mem[2445] = 4'b0000;
	mem[2446] = 4'b0000;
	mem[2447] = 4'b0000;
	mem[2448] = 4'b0000;
	mem[2449] = 4'b0000;
	mem[2450] = 4'b0000;
	mem[2451] = 4'b0000;
	mem[2452] = 4'b0000;
	mem[2453] = 4'b0000;
	mem[2454] = 4'b0000;
	mem[2455] = 4'b0000;
	mem[2456] = 4'b0000;
	mem[2457] = 4'b0001;
	mem[2458] = 4'b0001;
	mem[2459] = 4'b0000;
	mem[2460] = 4'b0000;
	mem[2461] = 4'b0000;
	mem[2462] = 4'b0000;
	mem[2463] = 4'b0000;
	mem[2464] = 4'b0000;
	mem[2465] = 4'b0000;
	mem[2466] = 4'b0000;
	mem[2467] = 4'b0000;
	mem[2468] = 4'b0000;
	mem[2469] = 4'b0000;
	mem[2470] = 4'b0000;
	mem[2471] = 4'b0000;
	mem[2472] = 4'b0000;
	mem[2473] = 4'b0000;
	mem[2474] = 4'b0000;
	mem[2475] = 4'b0000;
	mem[2476] = 4'b0000;
	mem[2477] = 4'b0000;
	mem[2478] = 4'b0000;
	mem[2479] = 4'b0000;
	mem[2480] = 4'b0000;
	mem[2481] = 4'b0000;
	mem[2482] = 4'b0000;
	mem[2483] = 4'b0000;
	mem[2484] = 4'b0000;
	mem[2485] = 4'b0000;
	mem[2486] = 4'b0000;
	mem[2487] = 4'b0000;
	mem[2488] = 4'b0000;
	mem[2489] = 4'b0000;
	mem[2490] = 4'b0000;
	mem[2491] = 4'b0000;
	mem[2492] = 4'b0000;
	mem[2493] = 4'b0000;
	mem[2494] = 4'b0000;
	mem[2495] = 4'b0000;
	mem[2496] = 4'b0000;
	mem[2497] = 4'b0000;
	mem[2498] = 4'b0000;
	mem[2499] = 4'b0000;
	mem[2500] = 4'b0001;
	mem[2501] = 4'b0000;
	mem[2502] = 4'b0000;
	mem[2503] = 4'b0000;
	mem[2504] = 4'b0000;
	mem[2505] = 4'b0000;
	mem[2506] = 4'b0000;
	mem[2507] = 4'b0000;
	mem[2508] = 4'b0000;
	mem[2509] = 4'b0000;
	mem[2510] = 4'b0000;
	mem[2511] = 4'b0000;
	mem[2512] = 4'b0000;
	mem[2513] = 4'b0000;
	mem[2514] = 4'b0000;
	mem[2515] = 4'b0000;
	mem[2516] = 4'b0000;
	mem[2517] = 4'b0000;
	mem[2518] = 4'b0000;
	mem[2519] = 4'b0000;
	mem[2520] = 4'b0000;
	mem[2521] = 4'b0000;
	mem[2522] = 4'b0000;
	mem[2523] = 4'b0000;
	mem[2524] = 4'b0000;
	mem[2525] = 4'b0000;
	mem[2526] = 4'b0000;
	mem[2527] = 4'b0000;
	mem[2528] = 4'b0000;
	mem[2529] = 4'b0000;
	mem[2530] = 4'b0000;
	mem[2531] = 4'b0000;
	mem[2532] = 4'b0000;
	mem[2533] = 4'b0000;
	mem[2534] = 4'b0000;
	mem[2535] = 4'b0000;
	mem[2536] = 4'b0000;
	mem[2537] = 4'b0000;
	mem[2538] = 4'b0000;
	mem[2539] = 4'b0000;
	mem[2540] = 4'b0000;
	mem[2541] = 4'b0000;
	mem[2542] = 4'b0000;
	mem[2543] = 4'b0000;
	mem[2544] = 4'b0000;
	mem[2545] = 4'b0000;
	mem[2546] = 4'b0000;
	mem[2547] = 4'b0000;
	mem[2548] = 4'b0000;
	mem[2549] = 4'b0000;
	mem[2550] = 4'b0000;
	mem[2551] = 4'b0000;
	mem[2552] = 4'b0000;
	mem[2553] = 4'b0000;
	mem[2554] = 4'b0000;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b0000;
	mem[2564] = 4'b0000;
	mem[2565] = 4'b0000;
	mem[2566] = 4'b0000;
	mem[2567] = 4'b0000;
	mem[2568] = 4'b0000;
	mem[2569] = 4'b0000;
	mem[2570] = 4'b0000;
	mem[2571] = 4'b0000;
	mem[2572] = 4'b0000;
	mem[2573] = 4'b0000;
	mem[2574] = 4'b0000;
	mem[2575] = 4'b0000;
	mem[2576] = 4'b0000;
	mem[2577] = 4'b0000;
	mem[2578] = 4'b0000;
	mem[2579] = 4'b0001;
	mem[2580] = 4'b0001;
	mem[2581] = 4'b0001;
	mem[2582] = 4'b0001;
	mem[2583] = 4'b0001;
	mem[2584] = 4'b0001;
	mem[2585] = 4'b0000;
	mem[2586] = 4'b0000;
	mem[2587] = 4'b0000;
	mem[2588] = 4'b0000;
	mem[2589] = 4'b0000;
	mem[2590] = 4'b0000;
	mem[2591] = 4'b0000;
	mem[2592] = 4'b0000;
	mem[2593] = 4'b0000;
	mem[2594] = 4'b0000;
	mem[2595] = 4'b0000;
	mem[2596] = 4'b0000;
	mem[2597] = 4'b0000;
	mem[2598] = 4'b0000;
	mem[2599] = 4'b0000;
	mem[2600] = 4'b0000;
	mem[2601] = 4'b0000;
	mem[2602] = 4'b0000;
	mem[2603] = 4'b0000;
	mem[2604] = 4'b0000;
	mem[2605] = 4'b0000;
	mem[2606] = 4'b0000;
	mem[2607] = 4'b0000;
	mem[2608] = 4'b0000;
	mem[2609] = 4'b0000;
	mem[2610] = 4'b0000;
	mem[2611] = 4'b0000;
	mem[2612] = 4'b0000;
	mem[2613] = 4'b0000;
	mem[2614] = 4'b0000;
	mem[2615] = 4'b0000;
	mem[2616] = 4'b0000;
	mem[2617] = 4'b0000;
	mem[2618] = 4'b0000;
	mem[2619] = 4'b0000;
	mem[2620] = 4'b0000;
	mem[2621] = 4'b0000;
	mem[2622] = 4'b0000;
	mem[2623] = 4'b0000;
	mem[2624] = 4'b0000;
	mem[2625] = 4'b0000;
	mem[2626] = 4'b0000;
	mem[2627] = 4'b0001;
	mem[2628] = 4'b0001;
	mem[2629] = 4'b0000;
	mem[2630] = 4'b0000;
	mem[2631] = 4'b0000;
	mem[2632] = 4'b0000;
	mem[2633] = 4'b0000;
	mem[2634] = 4'b0000;
	mem[2635] = 4'b0000;
	mem[2636] = 4'b0000;
	mem[2637] = 4'b0000;
	mem[2638] = 4'b0000;
	mem[2639] = 4'b0000;
	mem[2640] = 4'b0000;
	mem[2641] = 4'b0000;
	mem[2642] = 4'b0000;
	mem[2643] = 4'b0000;
	mem[2644] = 4'b0000;
	mem[2645] = 4'b0000;
	mem[2646] = 4'b0000;
	mem[2647] = 4'b0000;
	mem[2648] = 4'b0000;
	mem[2649] = 4'b0000;
	mem[2650] = 4'b0000;
	mem[2651] = 4'b0000;
	mem[2652] = 4'b0000;
	mem[2653] = 4'b0000;
	mem[2654] = 4'b0000;
	mem[2655] = 4'b0000;
	mem[2656] = 4'b0000;
	mem[2657] = 4'b0000;
	mem[2658] = 4'b0000;
	mem[2659] = 4'b0000;
	mem[2660] = 4'b0000;
	mem[2661] = 4'b0000;
	mem[2662] = 4'b0000;
	mem[2663] = 4'b0000;
	mem[2664] = 4'b0000;
	mem[2665] = 4'b0000;
	mem[2666] = 4'b0000;
	mem[2667] = 4'b0000;
	mem[2668] = 4'b0000;
	mem[2669] = 4'b0000;
	mem[2670] = 4'b0000;
	mem[2671] = 4'b0000;
	mem[2672] = 4'b0000;
	mem[2673] = 4'b0000;
	mem[2674] = 4'b0000;
	mem[2675] = 4'b0000;
	mem[2676] = 4'b0000;
	mem[2677] = 4'b0000;
	mem[2678] = 4'b0000;
	mem[2679] = 4'b0000;
	mem[2680] = 4'b0000;
	mem[2681] = 4'b0000;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b0000;
	mem[2692] = 4'b0000;
	mem[2693] = 4'b0000;
	mem[2694] = 4'b0000;
	mem[2695] = 4'b0000;
	mem[2696] = 4'b0000;
	mem[2697] = 4'b0000;
	mem[2698] = 4'b0000;
	mem[2699] = 4'b0000;
	mem[2700] = 4'b0000;
	mem[2701] = 4'b0000;
	mem[2702] = 4'b0000;
	mem[2703] = 4'b0000;
	mem[2704] = 4'b0000;
	mem[2705] = 4'b0000;
	mem[2706] = 4'b0000;
	mem[2707] = 4'b0000;
	mem[2708] = 4'b0000;
	mem[2709] = 4'b0000;
	mem[2710] = 4'b0000;
	mem[2711] = 4'b0000;
	mem[2712] = 4'b0000;
	mem[2713] = 4'b0000;
	mem[2714] = 4'b0000;
	mem[2715] = 4'b0000;
	mem[2716] = 4'b0000;
	mem[2717] = 4'b0000;
	mem[2718] = 4'b0000;
	mem[2719] = 4'b0000;
	mem[2720] = 4'b0000;
	mem[2721] = 4'b0000;
	mem[2722] = 4'b0000;
	mem[2723] = 4'b0000;
	mem[2724] = 4'b0000;
	mem[2725] = 4'b0000;
	mem[2726] = 4'b0000;
	mem[2727] = 4'b0000;
	mem[2728] = 4'b0000;
	mem[2729] = 4'b0000;
	mem[2730] = 4'b0000;
	mem[2731] = 4'b0000;
	mem[2732] = 4'b0000;
	mem[2733] = 4'b0000;
	mem[2734] = 4'b0000;
	mem[2735] = 4'b0000;
	mem[2736] = 4'b0000;
	mem[2737] = 4'b0000;
	mem[2738] = 4'b0000;
	mem[2739] = 4'b0000;
	mem[2740] = 4'b0000;
	mem[2741] = 4'b0000;
	mem[2742] = 4'b0000;
	mem[2743] = 4'b0000;
	mem[2744] = 4'b0000;
	mem[2745] = 4'b0000;
	mem[2746] = 4'b0000;
	mem[2747] = 4'b0000;
	mem[2748] = 4'b0000;
	mem[2749] = 4'b0000;
	mem[2750] = 4'b0001;
	mem[2751] = 4'b0000;
	mem[2752] = 4'b0000;
	mem[2753] = 4'b0000;
	mem[2754] = 4'b0001;
	mem[2755] = 4'b0001;
	mem[2756] = 4'b0000;
	mem[2757] = 4'b0000;
	mem[2758] = 4'b0000;
	mem[2759] = 4'b0000;
	mem[2760] = 4'b0000;
	mem[2761] = 4'b0000;
	mem[2762] = 4'b0000;
	mem[2763] = 4'b0000;
	mem[2764] = 4'b0000;
	mem[2765] = 4'b0000;
	mem[2766] = 4'b0000;
	mem[2767] = 4'b0000;
	mem[2768] = 4'b0000;
	mem[2769] = 4'b0000;
	mem[2770] = 4'b0000;
	mem[2771] = 4'b0000;
	mem[2772] = 4'b0000;
	mem[2773] = 4'b0000;
	mem[2774] = 4'b0000;
	mem[2775] = 4'b0000;
	mem[2776] = 4'b0000;
	mem[2777] = 4'b0000;
	mem[2778] = 4'b0000;
	mem[2779] = 4'b0000;
	mem[2780] = 4'b0000;
	mem[2781] = 4'b0000;
	mem[2782] = 4'b0000;
	mem[2783] = 4'b0000;
	mem[2784] = 4'b0000;
	mem[2785] = 4'b0000;
	mem[2786] = 4'b0000;
	mem[2787] = 4'b0000;
	mem[2788] = 4'b0000;
	mem[2789] = 4'b0000;
	mem[2790] = 4'b0000;
	mem[2791] = 4'b0000;
	mem[2792] = 4'b0000;
	mem[2793] = 4'b0000;
	mem[2794] = 4'b0000;
	mem[2795] = 4'b0000;
	mem[2796] = 4'b0000;
	mem[2797] = 4'b0000;
	mem[2798] = 4'b0000;
	mem[2799] = 4'b0000;
	mem[2800] = 4'b0000;
	mem[2801] = 4'b0000;
	mem[2802] = 4'b0000;
	mem[2803] = 4'b0000;
	mem[2804] = 4'b0000;
	mem[2805] = 4'b0000;
	mem[2806] = 4'b0000;
	mem[2807] = 4'b0000;
	mem[2808] = 4'b0000;
	mem[2809] = 4'b0000;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b0000;
	mem[2820] = 4'b0000;
	mem[2821] = 4'b0000;
	mem[2822] = 4'b0000;
	mem[2823] = 4'b0000;
	mem[2824] = 4'b0000;
	mem[2825] = 4'b0000;
	mem[2826] = 4'b0000;
	mem[2827] = 4'b0000;
	mem[2828] = 4'b0000;
	mem[2829] = 4'b0000;
	mem[2830] = 4'b0000;
	mem[2831] = 4'b0000;
	mem[2832] = 4'b0000;
	mem[2833] = 4'b0000;
	mem[2834] = 4'b0000;
	mem[2835] = 4'b0000;
	mem[2836] = 4'b0000;
	mem[2837] = 4'b0000;
	mem[2838] = 4'b0000;
	mem[2839] = 4'b0000;
	mem[2840] = 4'b0000;
	mem[2841] = 4'b0000;
	mem[2842] = 4'b0000;
	mem[2843] = 4'b0000;
	mem[2844] = 4'b0000;
	mem[2845] = 4'b0000;
	mem[2846] = 4'b0000;
	mem[2847] = 4'b0000;
	mem[2848] = 4'b0000;
	mem[2849] = 4'b0000;
	mem[2850] = 4'b0000;
	mem[2851] = 4'b0000;
	mem[2852] = 4'b0000;
	mem[2853] = 4'b0000;
	mem[2854] = 4'b0000;
	mem[2855] = 4'b0000;
	mem[2856] = 4'b0000;
	mem[2857] = 4'b0000;
	mem[2858] = 4'b0000;
	mem[2859] = 4'b0000;
	mem[2860] = 4'b0000;
	mem[2861] = 4'b0000;
	mem[2862] = 4'b0000;
	mem[2863] = 4'b0000;
	mem[2864] = 4'b0000;
	mem[2865] = 4'b0000;
	mem[2866] = 4'b0000;
	mem[2867] = 4'b0000;
	mem[2868] = 4'b0000;
	mem[2869] = 4'b0000;
	mem[2870] = 4'b0000;
	mem[2871] = 4'b0000;
	mem[2872] = 4'b0000;
	mem[2873] = 4'b0000;
	mem[2874] = 4'b0000;
	mem[2875] = 4'b0000;
	mem[2876] = 4'b0000;
	mem[2877] = 4'b0000;
	mem[2878] = 4'b0000;
	mem[2879] = 4'b0000;
	mem[2880] = 4'b0001;
	mem[2881] = 4'b0001;
	mem[2882] = 4'b0000;
	mem[2883] = 4'b0000;
	mem[2884] = 4'b0000;
	mem[2885] = 4'b0000;
	mem[2886] = 4'b0000;
	mem[2887] = 4'b0000;
	mem[2888] = 4'b0000;
	mem[2889] = 4'b0000;
	mem[2890] = 4'b0000;
	mem[2891] = 4'b0000;
	mem[2892] = 4'b0000;
	mem[2893] = 4'b0000;
	mem[2894] = 4'b0000;
	mem[2895] = 4'b0000;
	mem[2896] = 4'b0000;
	mem[2897] = 4'b0000;
	mem[2898] = 4'b0000;
	mem[2899] = 4'b0000;
	mem[2900] = 4'b0000;
	mem[2901] = 4'b0000;
	mem[2902] = 4'b0000;
	mem[2903] = 4'b0000;
	mem[2904] = 4'b0000;
	mem[2905] = 4'b0000;
	mem[2906] = 4'b0000;
	mem[2907] = 4'b0000;
	mem[2908] = 4'b0000;
	mem[2909] = 4'b0000;
	mem[2910] = 4'b0000;
	mem[2911] = 4'b0000;
	mem[2912] = 4'b0000;
	mem[2913] = 4'b0000;
	mem[2914] = 4'b0000;
	mem[2915] = 4'b0000;
	mem[2916] = 4'b0000;
	mem[2917] = 4'b0000;
	mem[2918] = 4'b0000;
	mem[2919] = 4'b0000;
	mem[2920] = 4'b0000;
	mem[2921] = 4'b0000;
	mem[2922] = 4'b0000;
	mem[2923] = 4'b0000;
	mem[2924] = 4'b0000;
	mem[2925] = 4'b0000;
	mem[2926] = 4'b0000;
	mem[2927] = 4'b0000;
	mem[2928] = 4'b0000;
	mem[2929] = 4'b0000;
	mem[2930] = 4'b0000;
	mem[2931] = 4'b0000;
	mem[2932] = 4'b0000;
	mem[2933] = 4'b0000;
	mem[2934] = 4'b0000;
	mem[2935] = 4'b0000;
	mem[2936] = 4'b0000;
	mem[2937] = 4'b0000;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b0000;
	mem[2948] = 4'b0000;
	mem[2949] = 4'b0000;
	mem[2950] = 4'b0000;
	mem[2951] = 4'b0000;
	mem[2952] = 4'b0000;
	mem[2953] = 4'b0000;
	mem[2954] = 4'b0000;
	mem[2955] = 4'b0000;
	mem[2956] = 4'b0000;
	mem[2957] = 4'b0000;
	mem[2958] = 4'b0000;
	mem[2959] = 4'b0000;
	mem[2960] = 4'b0000;
	mem[2961] = 4'b0000;
	mem[2962] = 4'b0000;
	mem[2963] = 4'b0000;
	mem[2964] = 4'b0000;
	mem[2965] = 4'b0000;
	mem[2966] = 4'b0000;
	mem[2967] = 4'b0000;
	mem[2968] = 4'b0000;
	mem[2969] = 4'b0000;
	mem[2970] = 4'b0000;
	mem[2971] = 4'b0000;
	mem[2972] = 4'b0000;
	mem[2973] = 4'b0000;
	mem[2974] = 4'b0000;
	mem[2975] = 4'b0000;
	mem[2976] = 4'b0000;
	mem[2977] = 4'b0000;
	mem[2978] = 4'b0000;
	mem[2979] = 4'b0000;
	mem[2980] = 4'b0000;
	mem[2981] = 4'b0000;
	mem[2982] = 4'b0000;
	mem[2983] = 4'b0000;
	mem[2984] = 4'b0000;
	mem[2985] = 4'b0000;
	mem[2986] = 4'b0000;
	mem[2987] = 4'b0000;
	mem[2988] = 4'b0000;
	mem[2989] = 4'b0000;
	mem[2990] = 4'b0000;
	mem[2991] = 4'b0000;
	mem[2992] = 4'b0000;
	mem[2993] = 4'b0000;
	mem[2994] = 4'b0000;
	mem[2995] = 4'b0000;
	mem[2996] = 4'b0000;
	mem[2997] = 4'b0000;
	mem[2998] = 4'b0000;
	mem[2999] = 4'b0000;
	mem[3000] = 4'b0000;
	mem[3001] = 4'b0000;
	mem[3002] = 4'b0000;
	mem[3003] = 4'b0000;
	mem[3004] = 4'b0000;
	mem[3005] = 4'b0000;
	mem[3006] = 4'b0000;
	mem[3007] = 4'b0000;
	mem[3008] = 4'b0000;
	mem[3009] = 4'b0000;
	mem[3010] = 4'b0000;
	mem[3011] = 4'b0000;
	mem[3012] = 4'b0000;
	mem[3013] = 4'b0000;
	mem[3014] = 4'b0000;
	mem[3015] = 4'b0000;
	mem[3016] = 4'b0000;
	mem[3017] = 4'b0000;
	mem[3018] = 4'b0000;
	mem[3019] = 4'b0000;
	mem[3020] = 4'b0000;
	mem[3021] = 4'b0000;
	mem[3022] = 4'b0000;
	mem[3023] = 4'b0000;
	mem[3024] = 4'b0000;
	mem[3025] = 4'b0000;
	mem[3026] = 4'b0000;
	mem[3027] = 4'b0000;
	mem[3028] = 4'b0000;
	mem[3029] = 4'b0000;
	mem[3030] = 4'b0000;
	mem[3031] = 4'b0000;
	mem[3032] = 4'b0000;
	mem[3033] = 4'b0000;
	mem[3034] = 4'b0000;
	mem[3035] = 4'b0000;
	mem[3036] = 4'b0000;
	mem[3037] = 4'b0000;
	mem[3038] = 4'b0000;
	mem[3039] = 4'b0000;
	mem[3040] = 4'b0000;
	mem[3041] = 4'b0000;
	mem[3042] = 4'b0000;
	mem[3043] = 4'b0000;
	mem[3044] = 4'b0000;
	mem[3045] = 4'b0000;
	mem[3046] = 4'b0000;
	mem[3047] = 4'b0000;
	mem[3048] = 4'b0000;
	mem[3049] = 4'b0000;
	mem[3050] = 4'b0000;
	mem[3051] = 4'b0000;
	mem[3052] = 4'b0000;
	mem[3053] = 4'b0000;
	mem[3054] = 4'b0000;
	mem[3055] = 4'b0000;
	mem[3056] = 4'b0000;
	mem[3057] = 4'b0000;
	mem[3058] = 4'b0000;
	mem[3059] = 4'b0000;
	mem[3060] = 4'b0000;
	mem[3061] = 4'b0000;
	mem[3062] = 4'b0000;
	mem[3063] = 4'b0000;
	mem[3064] = 4'b0000;
	mem[3065] = 4'b0000;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b0000;
	mem[3076] = 4'b0000;
	mem[3077] = 4'b0000;
	mem[3078] = 4'b0000;
	mem[3079] = 4'b0000;
	mem[3080] = 4'b0000;
	mem[3081] = 4'b0000;
	mem[3082] = 4'b0000;
	mem[3083] = 4'b0000;
	mem[3084] = 4'b0000;
	mem[3085] = 4'b0000;
	mem[3086] = 4'b0000;
	mem[3087] = 4'b0000;
	mem[3088] = 4'b0000;
	mem[3089] = 4'b0000;
	mem[3090] = 4'b0000;
	mem[3091] = 4'b0000;
	mem[3092] = 4'b0000;
	mem[3093] = 4'b0000;
	mem[3094] = 4'b0000;
	mem[3095] = 4'b0000;
	mem[3096] = 4'b0000;
	mem[3097] = 4'b0000;
	mem[3098] = 4'b0000;
	mem[3099] = 4'b0000;
	mem[3100] = 4'b0000;
	mem[3101] = 4'b0000;
	mem[3102] = 4'b0000;
	mem[3103] = 4'b0000;
	mem[3104] = 4'b0000;
	mem[3105] = 4'b0000;
	mem[3106] = 4'b0000;
	mem[3107] = 4'b0000;
	mem[3108] = 4'b0000;
	mem[3109] = 4'b0000;
	mem[3110] = 4'b0000;
	mem[3111] = 4'b0000;
	mem[3112] = 4'b0000;
	mem[3113] = 4'b0000;
	mem[3114] = 4'b0000;
	mem[3115] = 4'b0000;
	mem[3116] = 4'b0000;
	mem[3117] = 4'b0000;
	mem[3118] = 4'b0000;
	mem[3119] = 4'b0000;
	mem[3120] = 4'b0000;
	mem[3121] = 4'b0000;
	mem[3122] = 4'b0000;
	mem[3123] = 4'b0000;
	mem[3124] = 4'b0000;
	mem[3125] = 4'b0000;
	mem[3126] = 4'b0000;
	mem[3127] = 4'b0000;
	mem[3128] = 4'b0000;
	mem[3129] = 4'b0000;
	mem[3130] = 4'b0000;
	mem[3131] = 4'b0000;
	mem[3132] = 4'b0000;
	mem[3133] = 4'b0000;
	mem[3134] = 4'b0000;
	mem[3135] = 4'b0000;
	mem[3136] = 4'b0000;
	mem[3137] = 4'b0000;
	mem[3138] = 4'b0000;
	mem[3139] = 4'b0000;
	mem[3140] = 4'b0000;
	mem[3141] = 4'b0000;
	mem[3142] = 4'b0000;
	mem[3143] = 4'b0000;
	mem[3144] = 4'b0000;
	mem[3145] = 4'b0000;
	mem[3146] = 4'b0000;
	mem[3147] = 4'b0000;
	mem[3148] = 4'b0000;
	mem[3149] = 4'b0000;
	mem[3150] = 4'b0000;
	mem[3151] = 4'b0000;
	mem[3152] = 4'b0000;
	mem[3153] = 4'b0000;
	mem[3154] = 4'b0000;
	mem[3155] = 4'b0000;
	mem[3156] = 4'b0000;
	mem[3157] = 4'b0000;
	mem[3158] = 4'b0000;
	mem[3159] = 4'b0000;
	mem[3160] = 4'b0000;
	mem[3161] = 4'b0000;
	mem[3162] = 4'b0000;
	mem[3163] = 4'b0000;
	mem[3164] = 4'b0000;
	mem[3165] = 4'b0000;
	mem[3166] = 4'b0000;
	mem[3167] = 4'b0000;
	mem[3168] = 4'b0000;
	mem[3169] = 4'b0000;
	mem[3170] = 4'b0000;
	mem[3171] = 4'b0000;
	mem[3172] = 4'b0000;
	mem[3173] = 4'b0000;
	mem[3174] = 4'b0000;
	mem[3175] = 4'b0000;
	mem[3176] = 4'b0000;
	mem[3177] = 4'b0000;
	mem[3178] = 4'b0000;
	mem[3179] = 4'b0000;
	mem[3180] = 4'b0000;
	mem[3181] = 4'b0000;
	mem[3182] = 4'b0000;
	mem[3183] = 4'b0000;
	mem[3184] = 4'b0000;
	mem[3185] = 4'b0000;
	mem[3186] = 4'b0000;
	mem[3187] = 4'b0000;
	mem[3188] = 4'b0000;
	mem[3189] = 4'b0000;
	mem[3190] = 4'b0000;
	mem[3191] = 4'b0000;
	mem[3192] = 4'b0000;
	mem[3193] = 4'b0000;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b0000;
	mem[3204] = 4'b0000;
	mem[3205] = 4'b0000;
	mem[3206] = 4'b0000;
	mem[3207] = 4'b0000;
	mem[3208] = 4'b0000;
	mem[3209] = 4'b0000;
	mem[3210] = 4'b0000;
	mem[3211] = 4'b0000;
	mem[3212] = 4'b0000;
	mem[3213] = 4'b0000;
	mem[3214] = 4'b0000;
	mem[3215] = 4'b0000;
	mem[3216] = 4'b0000;
	mem[3217] = 4'b0000;
	mem[3218] = 4'b0000;
	mem[3219] = 4'b0000;
	mem[3220] = 4'b0000;
	mem[3221] = 4'b0000;
	mem[3222] = 4'b0000;
	mem[3223] = 4'b0000;
	mem[3224] = 4'b0000;
	mem[3225] = 4'b0000;
	mem[3226] = 4'b0000;
	mem[3227] = 4'b0000;
	mem[3228] = 4'b0000;
	mem[3229] = 4'b0000;
	mem[3230] = 4'b0000;
	mem[3231] = 4'b0000;
	mem[3232] = 4'b0000;
	mem[3233] = 4'b0000;
	mem[3234] = 4'b0000;
	mem[3235] = 4'b0000;
	mem[3236] = 4'b0000;
	mem[3237] = 4'b0000;
	mem[3238] = 4'b0000;
	mem[3239] = 4'b0000;
	mem[3240] = 4'b0000;
	mem[3241] = 4'b0000;
	mem[3242] = 4'b0000;
	mem[3243] = 4'b0000;
	mem[3244] = 4'b0000;
	mem[3245] = 4'b0000;
	mem[3246] = 4'b0000;
	mem[3247] = 4'b0000;
	mem[3248] = 4'b0000;
	mem[3249] = 4'b0000;
	mem[3250] = 4'b0000;
	mem[3251] = 4'b0000;
	mem[3252] = 4'b0000;
	mem[3253] = 4'b0000;
	mem[3254] = 4'b0000;
	mem[3255] = 4'b0000;
	mem[3256] = 4'b0000;
	mem[3257] = 4'b0000;
	mem[3258] = 4'b0000;
	mem[3259] = 4'b0000;
	mem[3260] = 4'b0000;
	mem[3261] = 4'b0000;
	mem[3262] = 4'b0001;
	mem[3263] = 4'b0000;
	mem[3264] = 4'b0000;
	mem[3265] = 4'b0000;
	mem[3266] = 4'b0000;
	mem[3267] = 4'b0000;
	mem[3268] = 4'b0000;
	mem[3269] = 4'b0000;
	mem[3270] = 4'b0000;
	mem[3271] = 4'b0000;
	mem[3272] = 4'b0000;
	mem[3273] = 4'b0000;
	mem[3274] = 4'b0000;
	mem[3275] = 4'b0000;
	mem[3276] = 4'b0000;
	mem[3277] = 4'b0000;
	mem[3278] = 4'b0000;
	mem[3279] = 4'b0000;
	mem[3280] = 4'b0000;
	mem[3281] = 4'b0000;
	mem[3282] = 4'b0000;
	mem[3283] = 4'b0000;
	mem[3284] = 4'b0000;
	mem[3285] = 4'b0000;
	mem[3286] = 4'b0000;
	mem[3287] = 4'b0000;
	mem[3288] = 4'b0000;
	mem[3289] = 4'b0000;
	mem[3290] = 4'b0000;
	mem[3291] = 4'b0000;
	mem[3292] = 4'b0000;
	mem[3293] = 4'b0000;
	mem[3294] = 4'b0000;
	mem[3295] = 4'b0000;
	mem[3296] = 4'b0000;
	mem[3297] = 4'b0000;
	mem[3298] = 4'b0000;
	mem[3299] = 4'b0000;
	mem[3300] = 4'b0000;
	mem[3301] = 4'b0000;
	mem[3302] = 4'b0000;
	mem[3303] = 4'b0000;
	mem[3304] = 4'b0000;
	mem[3305] = 4'b0000;
	mem[3306] = 4'b0000;
	mem[3307] = 4'b0000;
	mem[3308] = 4'b0000;
	mem[3309] = 4'b0000;
	mem[3310] = 4'b0000;
	mem[3311] = 4'b0000;
	mem[3312] = 4'b0000;
	mem[3313] = 4'b0000;
	mem[3314] = 4'b0000;
	mem[3315] = 4'b0000;
	mem[3316] = 4'b0000;
	mem[3317] = 4'b0000;
	mem[3318] = 4'b0000;
	mem[3319] = 4'b0000;
	mem[3320] = 4'b0000;
	mem[3321] = 4'b0000;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b0000;
	mem[3332] = 4'b0000;
	mem[3333] = 4'b0000;
	mem[3334] = 4'b0000;
	mem[3335] = 4'b0000;
	mem[3336] = 4'b0000;
	mem[3337] = 4'b0000;
	mem[3338] = 4'b0000;
	mem[3339] = 4'b0000;
	mem[3340] = 4'b0000;
	mem[3341] = 4'b0000;
	mem[3342] = 4'b0000;
	mem[3343] = 4'b0000;
	mem[3344] = 4'b0000;
	mem[3345] = 4'b0000;
	mem[3346] = 4'b0001;
	mem[3347] = 4'b0001;
	mem[3348] = 4'b0000;
	mem[3349] = 4'b0000;
	mem[3350] = 4'b0000;
	mem[3351] = 4'b0000;
	mem[3352] = 4'b0000;
	mem[3353] = 4'b0000;
	mem[3354] = 4'b0000;
	mem[3355] = 4'b0000;
	mem[3356] = 4'b0000;
	mem[3357] = 4'b0000;
	mem[3358] = 4'b0000;
	mem[3359] = 4'b0000;
	mem[3360] = 4'b0000;
	mem[3361] = 4'b0000;
	mem[3362] = 4'b0000;
	mem[3363] = 4'b0000;
	mem[3364] = 4'b0000;
	mem[3365] = 4'b0000;
	mem[3366] = 4'b0000;
	mem[3367] = 4'b0000;
	mem[3368] = 4'b0000;
	mem[3369] = 4'b0000;
	mem[3370] = 4'b0000;
	mem[3371] = 4'b0000;
	mem[3372] = 4'b0000;
	mem[3373] = 4'b0000;
	mem[3374] = 4'b0000;
	mem[3375] = 4'b0000;
	mem[3376] = 4'b0000;
	mem[3377] = 4'b0000;
	mem[3378] = 4'b0000;
	mem[3379] = 4'b0000;
	mem[3380] = 4'b0000;
	mem[3381] = 4'b0000;
	mem[3382] = 4'b0000;
	mem[3383] = 4'b0000;
	mem[3384] = 4'b0000;
	mem[3385] = 4'b0000;
	mem[3386] = 4'b0000;
	mem[3387] = 4'b0000;
	mem[3388] = 4'b0000;
	mem[3389] = 4'b0001;
	mem[3390] = 4'b0001;
	mem[3391] = 4'b0000;
	mem[3392] = 4'b0000;
	mem[3393] = 4'b0000;
	mem[3394] = 4'b0000;
	mem[3395] = 4'b0000;
	mem[3396] = 4'b0000;
	mem[3397] = 4'b0000;
	mem[3398] = 4'b0000;
	mem[3399] = 4'b0000;
	mem[3400] = 4'b0000;
	mem[3401] = 4'b0000;
	mem[3402] = 4'b0000;
	mem[3403] = 4'b0000;
	mem[3404] = 4'b0000;
	mem[3405] = 4'b0000;
	mem[3406] = 4'b0000;
	mem[3407] = 4'b0000;
	mem[3408] = 4'b0000;
	mem[3409] = 4'b0000;
	mem[3410] = 4'b0000;
	mem[3411] = 4'b0000;
	mem[3412] = 4'b0000;
	mem[3413] = 4'b0000;
	mem[3414] = 4'b0000;
	mem[3415] = 4'b0000;
	mem[3416] = 4'b0000;
	mem[3417] = 4'b0000;
	mem[3418] = 4'b0000;
	mem[3419] = 4'b0000;
	mem[3420] = 4'b0000;
	mem[3421] = 4'b0000;
	mem[3422] = 4'b0000;
	mem[3423] = 4'b0000;
	mem[3424] = 4'b0000;
	mem[3425] = 4'b0000;
	mem[3426] = 4'b0000;
	mem[3427] = 4'b0000;
	mem[3428] = 4'b0000;
	mem[3429] = 4'b0000;
	mem[3430] = 4'b0000;
	mem[3431] = 4'b0000;
	mem[3432] = 4'b0000;
	mem[3433] = 4'b0000;
	mem[3434] = 4'b0000;
	mem[3435] = 4'b0000;
	mem[3436] = 4'b0000;
	mem[3437] = 4'b0000;
	mem[3438] = 4'b0000;
	mem[3439] = 4'b0000;
	mem[3440] = 4'b0000;
	mem[3441] = 4'b0000;
	mem[3442] = 4'b0000;
	mem[3443] = 4'b0000;
	mem[3444] = 4'b0000;
	mem[3445] = 4'b0000;
	mem[3446] = 4'b0000;
	mem[3447] = 4'b0000;
	mem[3448] = 4'b0000;
	mem[3449] = 4'b0000;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b0000;
	mem[3460] = 4'b0000;
	mem[3461] = 4'b0000;
	mem[3462] = 4'b0000;
	mem[3463] = 4'b0000;
	mem[3464] = 4'b0000;
	mem[3465] = 4'b0000;
	mem[3466] = 4'b0000;
	mem[3467] = 4'b0000;
	mem[3468] = 4'b0000;
	mem[3469] = 4'b0000;
	mem[3470] = 4'b0000;
	mem[3471] = 4'b0000;
	mem[3472] = 4'b0000;
	mem[3473] = 4'b0001;
	mem[3474] = 4'b0001;
	mem[3475] = 4'b0000;
	mem[3476] = 4'b0000;
	mem[3477] = 4'b0000;
	mem[3478] = 4'b0000;
	mem[3479] = 4'b0000;
	mem[3480] = 4'b0000;
	mem[3481] = 4'b0000;
	mem[3482] = 4'b0000;
	mem[3483] = 4'b0000;
	mem[3484] = 4'b0000;
	mem[3485] = 4'b0000;
	mem[3486] = 4'b0000;
	mem[3487] = 4'b0000;
	mem[3488] = 4'b0000;
	mem[3489] = 4'b0000;
	mem[3490] = 4'b0000;
	mem[3491] = 4'b0000;
	mem[3492] = 4'b0000;
	mem[3493] = 4'b0000;
	mem[3494] = 4'b0000;
	mem[3495] = 4'b0000;
	mem[3496] = 4'b0000;
	mem[3497] = 4'b0000;
	mem[3498] = 4'b0000;
	mem[3499] = 4'b0000;
	mem[3500] = 4'b0000;
	mem[3501] = 4'b0000;
	mem[3502] = 4'b0000;
	mem[3503] = 4'b0000;
	mem[3504] = 4'b0000;
	mem[3505] = 4'b0000;
	mem[3506] = 4'b0000;
	mem[3507] = 4'b0000;
	mem[3508] = 4'b0000;
	mem[3509] = 4'b0000;
	mem[3510] = 4'b0000;
	mem[3511] = 4'b0000;
	mem[3512] = 4'b0000;
	mem[3513] = 4'b0000;
	mem[3514] = 4'b0000;
	mem[3515] = 4'b0000;
	mem[3516] = 4'b0000;
	mem[3517] = 4'b0000;
	mem[3518] = 4'b0000;
	mem[3519] = 4'b0000;
	mem[3520] = 4'b0000;
	mem[3521] = 4'b0000;
	mem[3522] = 4'b0000;
	mem[3523] = 4'b0000;
	mem[3524] = 4'b0000;
	mem[3525] = 4'b0000;
	mem[3526] = 4'b0000;
	mem[3527] = 4'b0000;
	mem[3528] = 4'b0000;
	mem[3529] = 4'b0000;
	mem[3530] = 4'b0000;
	mem[3531] = 4'b0000;
	mem[3532] = 4'b0000;
	mem[3533] = 4'b0000;
	mem[3534] = 4'b0000;
	mem[3535] = 4'b0000;
	mem[3536] = 4'b0000;
	mem[3537] = 4'b0000;
	mem[3538] = 4'b0000;
	mem[3539] = 4'b0000;
	mem[3540] = 4'b0000;
	mem[3541] = 4'b0000;
	mem[3542] = 4'b0000;
	mem[3543] = 4'b0000;
	mem[3544] = 4'b0000;
	mem[3545] = 4'b0000;
	mem[3546] = 4'b0000;
	mem[3547] = 4'b0000;
	mem[3548] = 4'b0000;
	mem[3549] = 4'b0000;
	mem[3550] = 4'b0000;
	mem[3551] = 4'b0000;
	mem[3552] = 4'b0000;
	mem[3553] = 4'b0000;
	mem[3554] = 4'b0000;
	mem[3555] = 4'b0000;
	mem[3556] = 4'b0000;
	mem[3557] = 4'b0000;
	mem[3558] = 4'b0000;
	mem[3559] = 4'b0000;
	mem[3560] = 4'b0000;
	mem[3561] = 4'b0000;
	mem[3562] = 4'b0000;
	mem[3563] = 4'b0000;
	mem[3564] = 4'b0000;
	mem[3565] = 4'b0000;
	mem[3566] = 4'b0000;
	mem[3567] = 4'b0000;
	mem[3568] = 4'b0000;
	mem[3569] = 4'b0000;
	mem[3570] = 4'b0000;
	mem[3571] = 4'b0000;
	mem[3572] = 4'b0000;
	mem[3573] = 4'b0000;
	mem[3574] = 4'b0000;
	mem[3575] = 4'b0000;
	mem[3576] = 4'b0000;
	mem[3577] = 4'b0000;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b0000;
	mem[3588] = 4'b0000;
	mem[3589] = 4'b0000;
	mem[3590] = 4'b0000;
	mem[3591] = 4'b0000;
	mem[3592] = 4'b0000;
	mem[3593] = 4'b0000;
	mem[3594] = 4'b0000;
	mem[3595] = 4'b0000;
	mem[3596] = 4'b0000;
	mem[3597] = 4'b0000;
	mem[3598] = 4'b0000;
	mem[3599] = 4'b0000;
	mem[3600] = 4'b0001;
	mem[3601] = 4'b0001;
	mem[3602] = 4'b0000;
	mem[3603] = 4'b0000;
	mem[3604] = 4'b0000;
	mem[3605] = 4'b0000;
	mem[3606] = 4'b0000;
	mem[3607] = 4'b0000;
	mem[3608] = 4'b0000;
	mem[3609] = 4'b0000;
	mem[3610] = 4'b0000;
	mem[3611] = 4'b0000;
	mem[3612] = 4'b0000;
	mem[3613] = 4'b0000;
	mem[3614] = 4'b0000;
	mem[3615] = 4'b0000;
	mem[3616] = 4'b0000;
	mem[3617] = 4'b0000;
	mem[3618] = 4'b0000;
	mem[3619] = 4'b0000;
	mem[3620] = 4'b0000;
	mem[3621] = 4'b0000;
	mem[3622] = 4'b0000;
	mem[3623] = 4'b0000;
	mem[3624] = 4'b0000;
	mem[3625] = 4'b0000;
	mem[3626] = 4'b0000;
	mem[3627] = 4'b0000;
	mem[3628] = 4'b0000;
	mem[3629] = 4'b0000;
	mem[3630] = 4'b0000;
	mem[3631] = 4'b0000;
	mem[3632] = 4'b0000;
	mem[3633] = 4'b0000;
	mem[3634] = 4'b0000;
	mem[3635] = 4'b0000;
	mem[3636] = 4'b0000;
	mem[3637] = 4'b0000;
	mem[3638] = 4'b0000;
	mem[3639] = 4'b0000;
	mem[3640] = 4'b0000;
	mem[3641] = 4'b0000;
	mem[3642] = 4'b0000;
	mem[3643] = 4'b0000;
	mem[3644] = 4'b0000;
	mem[3645] = 4'b0000;
	mem[3646] = 4'b0000;
	mem[3647] = 4'b0000;
	mem[3648] = 4'b0000;
	mem[3649] = 4'b0000;
	mem[3650] = 4'b0000;
	mem[3651] = 4'b0000;
	mem[3652] = 4'b0000;
	mem[3653] = 4'b0000;
	mem[3654] = 4'b0000;
	mem[3655] = 4'b0000;
	mem[3656] = 4'b0000;
	mem[3657] = 4'b0000;
	mem[3658] = 4'b0000;
	mem[3659] = 4'b0000;
	mem[3660] = 4'b0000;
	mem[3661] = 4'b0000;
	mem[3662] = 4'b0000;
	mem[3663] = 4'b0000;
	mem[3664] = 4'b0000;
	mem[3665] = 4'b0000;
	mem[3666] = 4'b0000;
	mem[3667] = 4'b0000;
	mem[3668] = 4'b0000;
	mem[3669] = 4'b0000;
	mem[3670] = 4'b0000;
	mem[3671] = 4'b0000;
	mem[3672] = 4'b0000;
	mem[3673] = 4'b0000;
	mem[3674] = 4'b0000;
	mem[3675] = 4'b0000;
	mem[3676] = 4'b0000;
	mem[3677] = 4'b0000;
	mem[3678] = 4'b0000;
	mem[3679] = 4'b0000;
	mem[3680] = 4'b0000;
	mem[3681] = 4'b0000;
	mem[3682] = 4'b0000;
	mem[3683] = 4'b0000;
	mem[3684] = 4'b0000;
	mem[3685] = 4'b0000;
	mem[3686] = 4'b0000;
	mem[3687] = 4'b0000;
	mem[3688] = 4'b0000;
	mem[3689] = 4'b0000;
	mem[3690] = 4'b0000;
	mem[3691] = 4'b0000;
	mem[3692] = 4'b0000;
	mem[3693] = 4'b0000;
	mem[3694] = 4'b0000;
	mem[3695] = 4'b0000;
	mem[3696] = 4'b0000;
	mem[3697] = 4'b0000;
	mem[3698] = 4'b0000;
	mem[3699] = 4'b0000;
	mem[3700] = 4'b0000;
	mem[3701] = 4'b0000;
	mem[3702] = 4'b0000;
	mem[3703] = 4'b0000;
	mem[3704] = 4'b0000;
	mem[3705] = 4'b0000;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b0000;
	mem[3716] = 4'b0000;
	mem[3717] = 4'b0000;
	mem[3718] = 4'b0000;
	mem[3719] = 4'b0000;
	mem[3720] = 4'b0000;
	mem[3721] = 4'b0000;
	mem[3722] = 4'b0000;
	mem[3723] = 4'b0000;
	mem[3724] = 4'b0000;
	mem[3725] = 4'b0000;
	mem[3726] = 4'b0000;
	mem[3727] = 4'b0000;
	mem[3728] = 4'b0000;
	mem[3729] = 4'b0000;
	mem[3730] = 4'b0000;
	mem[3731] = 4'b0000;
	mem[3732] = 4'b0000;
	mem[3733] = 4'b0000;
	mem[3734] = 4'b0000;
	mem[3735] = 4'b0000;
	mem[3736] = 4'b0000;
	mem[3737] = 4'b0000;
	mem[3738] = 4'b0000;
	mem[3739] = 4'b0000;
	mem[3740] = 4'b0000;
	mem[3741] = 4'b0000;
	mem[3742] = 4'b0000;
	mem[3743] = 4'b0000;
	mem[3744] = 4'b0000;
	mem[3745] = 4'b0000;
	mem[3746] = 4'b0000;
	mem[3747] = 4'b0000;
	mem[3748] = 4'b0000;
	mem[3749] = 4'b0000;
	mem[3750] = 4'b0000;
	mem[3751] = 4'b0000;
	mem[3752] = 4'b0000;
	mem[3753] = 4'b0000;
	mem[3754] = 4'b0000;
	mem[3755] = 4'b0000;
	mem[3756] = 4'b0000;
	mem[3757] = 4'b0000;
	mem[3758] = 4'b0000;
	mem[3759] = 4'b0000;
	mem[3760] = 4'b0000;
	mem[3761] = 4'b0000;
	mem[3762] = 4'b0000;
	mem[3763] = 4'b0000;
	mem[3764] = 4'b0000;
	mem[3765] = 4'b0000;
	mem[3766] = 4'b0000;
	mem[3767] = 4'b0000;
	mem[3768] = 4'b0000;
	mem[3769] = 4'b0000;
	mem[3770] = 4'b0000;
	mem[3771] = 4'b0000;
	mem[3772] = 4'b0000;
	mem[3773] = 4'b0000;
	mem[3774] = 4'b0000;
	mem[3775] = 4'b0000;
	mem[3776] = 4'b0000;
	mem[3777] = 4'b0000;
	mem[3778] = 4'b0000;
	mem[3779] = 4'b0000;
	mem[3780] = 4'b0000;
	mem[3781] = 4'b0000;
	mem[3782] = 4'b0000;
	mem[3783] = 4'b0000;
	mem[3784] = 4'b0000;
	mem[3785] = 4'b0000;
	mem[3786] = 4'b0000;
	mem[3787] = 4'b0000;
	mem[3788] = 4'b0000;
	mem[3789] = 4'b0000;
	mem[3790] = 4'b0000;
	mem[3791] = 4'b0000;
	mem[3792] = 4'b0000;
	mem[3793] = 4'b0000;
	mem[3794] = 4'b0000;
	mem[3795] = 4'b0000;
	mem[3796] = 4'b0000;
	mem[3797] = 4'b0000;
	mem[3798] = 4'b0000;
	mem[3799] = 4'b0000;
	mem[3800] = 4'b0000;
	mem[3801] = 4'b0000;
	mem[3802] = 4'b0000;
	mem[3803] = 4'b0000;
	mem[3804] = 4'b0000;
	mem[3805] = 4'b0000;
	mem[3806] = 4'b0000;
	mem[3807] = 4'b0000;
	mem[3808] = 4'b0000;
	mem[3809] = 4'b0000;
	mem[3810] = 4'b0000;
	mem[3811] = 4'b0000;
	mem[3812] = 4'b0000;
	mem[3813] = 4'b0000;
	mem[3814] = 4'b0000;
	mem[3815] = 4'b0000;
	mem[3816] = 4'b0000;
	mem[3817] = 4'b0000;
	mem[3818] = 4'b0000;
	mem[3819] = 4'b0000;
	mem[3820] = 4'b0000;
	mem[3821] = 4'b0000;
	mem[3822] = 4'b0000;
	mem[3823] = 4'b0000;
	mem[3824] = 4'b0000;
	mem[3825] = 4'b0000;
	mem[3826] = 4'b0000;
	mem[3827] = 4'b0000;
	mem[3828] = 4'b0000;
	mem[3829] = 4'b0000;
	mem[3830] = 4'b0000;
	mem[3831] = 4'b0000;
	mem[3832] = 4'b0000;
	mem[3833] = 4'b0000;
	mem[3834] = 4'b0000;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b0000;
	mem[3844] = 4'b0000;
	mem[3845] = 4'b0000;
	mem[3846] = 4'b0000;
	mem[3847] = 4'b0000;
	mem[3848] = 4'b0000;
	mem[3849] = 4'b0000;
	mem[3850] = 4'b0000;
	mem[3851] = 4'b0000;
	mem[3852] = 4'b0000;
	mem[3853] = 4'b0000;
	mem[3854] = 4'b0000;
	mem[3855] = 4'b0000;
	mem[3856] = 4'b0000;
	mem[3857] = 4'b0000;
	mem[3858] = 4'b0000;
	mem[3859] = 4'b0000;
	mem[3860] = 4'b0000;
	mem[3861] = 4'b0000;
	mem[3862] = 4'b0000;
	mem[3863] = 4'b0000;
	mem[3864] = 4'b0000;
	mem[3865] = 4'b0000;
	mem[3866] = 4'b0000;
	mem[3867] = 4'b0000;
	mem[3868] = 4'b0000;
	mem[3869] = 4'b0000;
	mem[3870] = 4'b0000;
	mem[3871] = 4'b0000;
	mem[3872] = 4'b0000;
	mem[3873] = 4'b0000;
	mem[3874] = 4'b0000;
	mem[3875] = 4'b0000;
	mem[3876] = 4'b0000;
	mem[3877] = 4'b0000;
	mem[3878] = 4'b0000;
	mem[3879] = 4'b0000;
	mem[3880] = 4'b0000;
	mem[3881] = 4'b0000;
	mem[3882] = 4'b0000;
	mem[3883] = 4'b0000;
	mem[3884] = 4'b0000;
	mem[3885] = 4'b0000;
	mem[3886] = 4'b0000;
	mem[3887] = 4'b0000;
	mem[3888] = 4'b0000;
	mem[3889] = 4'b0000;
	mem[3890] = 4'b0000;
	mem[3891] = 4'b0000;
	mem[3892] = 4'b0000;
	mem[3893] = 4'b0000;
	mem[3894] = 4'b0000;
	mem[3895] = 4'b0000;
	mem[3896] = 4'b0000;
	mem[3897] = 4'b0000;
	mem[3898] = 4'b0000;
	mem[3899] = 4'b0000;
	mem[3900] = 4'b0000;
	mem[3901] = 4'b0000;
	mem[3902] = 4'b0000;
	mem[3903] = 4'b0000;
	mem[3904] = 4'b0000;
	mem[3905] = 4'b0000;
	mem[3906] = 4'b0000;
	mem[3907] = 4'b0000;
	mem[3908] = 4'b0000;
	mem[3909] = 4'b0000;
	mem[3910] = 4'b0000;
	mem[3911] = 4'b0000;
	mem[3912] = 4'b0000;
	mem[3913] = 4'b0000;
	mem[3914] = 4'b0000;
	mem[3915] = 4'b0000;
	mem[3916] = 4'b0000;
	mem[3917] = 4'b0000;
	mem[3918] = 4'b0000;
	mem[3919] = 4'b0000;
	mem[3920] = 4'b0000;
	mem[3921] = 4'b0000;
	mem[3922] = 4'b0000;
	mem[3923] = 4'b0000;
	mem[3924] = 4'b0000;
	mem[3925] = 4'b0000;
	mem[3926] = 4'b0000;
	mem[3927] = 4'b0000;
	mem[3928] = 4'b0000;
	mem[3929] = 4'b0000;
	mem[3930] = 4'b0000;
	mem[3931] = 4'b0000;
	mem[3932] = 4'b0000;
	mem[3933] = 4'b0000;
	mem[3934] = 4'b0000;
	mem[3935] = 4'b0000;
	mem[3936] = 4'b0000;
	mem[3937] = 4'b0000;
	mem[3938] = 4'b0000;
	mem[3939] = 4'b0000;
	mem[3940] = 4'b0000;
	mem[3941] = 4'b0000;
	mem[3942] = 4'b0000;
	mem[3943] = 4'b0000;
	mem[3944] = 4'b0000;
	mem[3945] = 4'b0000;
	mem[3946] = 4'b0000;
	mem[3947] = 4'b0000;
	mem[3948] = 4'b0000;
	mem[3949] = 4'b0000;
	mem[3950] = 4'b0000;
	mem[3951] = 4'b0000;
	mem[3952] = 4'b0000;
	mem[3953] = 4'b0000;
	mem[3954] = 4'b0000;
	mem[3955] = 4'b0000;
	mem[3956] = 4'b0000;
	mem[3957] = 4'b0000;
	mem[3958] = 4'b0000;
	mem[3959] = 4'b0000;
	mem[3960] = 4'b0000;
	mem[3961] = 4'b0000;
	mem[3962] = 4'b0000;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b0000;
	mem[3972] = 4'b0000;
	mem[3973] = 4'b0000;
	mem[3974] = 4'b0000;
	mem[3975] = 4'b0000;
	mem[3976] = 4'b0000;
	mem[3977] = 4'b0000;
	mem[3978] = 4'b0000;
	mem[3979] = 4'b0000;
	mem[3980] = 4'b0000;
	mem[3981] = 4'b0000;
	mem[3982] = 4'b0000;
	mem[3983] = 4'b0000;
	mem[3984] = 4'b0000;
	mem[3985] = 4'b0000;
	mem[3986] = 4'b0000;
	mem[3987] = 4'b0000;
	mem[3988] = 4'b0000;
	mem[3989] = 4'b0000;
	mem[3990] = 4'b0000;
	mem[3991] = 4'b0000;
	mem[3992] = 4'b0000;
	mem[3993] = 4'b0000;
	mem[3994] = 4'b0000;
	mem[3995] = 4'b0000;
	mem[3996] = 4'b0000;
	mem[3997] = 4'b0000;
	mem[3998] = 4'b0000;
	mem[3999] = 4'b0000;
	mem[4000] = 4'b0000;
	mem[4001] = 4'b0000;
	mem[4002] = 4'b0000;
	mem[4003] = 4'b0000;
	mem[4004] = 4'b0000;
	mem[4005] = 4'b0000;
	mem[4006] = 4'b0000;
	mem[4007] = 4'b0000;
	mem[4008] = 4'b0000;
	mem[4009] = 4'b0000;
	mem[4010] = 4'b0000;
	mem[4011] = 4'b0000;
	mem[4012] = 4'b0000;
	mem[4013] = 4'b0000;
	mem[4014] = 4'b0000;
	mem[4015] = 4'b0000;
	mem[4016] = 4'b0000;
	mem[4017] = 4'b0000;
	mem[4018] = 4'b0000;
	mem[4019] = 4'b0000;
	mem[4020] = 4'b0000;
	mem[4021] = 4'b0000;
	mem[4022] = 4'b0000;
	mem[4023] = 4'b0000;
	mem[4024] = 4'b0000;
	mem[4025] = 4'b0000;
	mem[4026] = 4'b0000;
	mem[4027] = 4'b0000;
	mem[4028] = 4'b0000;
	mem[4029] = 4'b0000;
	mem[4030] = 4'b0000;
	mem[4031] = 4'b0000;
	mem[4032] = 4'b0000;
	mem[4033] = 4'b0000;
	mem[4034] = 4'b0000;
	mem[4035] = 4'b0000;
	mem[4036] = 4'b0000;
	mem[4037] = 4'b0000;
	mem[4038] = 4'b0000;
	mem[4039] = 4'b0000;
	mem[4040] = 4'b0000;
	mem[4041] = 4'b0000;
	mem[4042] = 4'b0000;
	mem[4043] = 4'b0000;
	mem[4044] = 4'b0000;
	mem[4045] = 4'b0000;
	mem[4046] = 4'b0000;
	mem[4047] = 4'b0000;
	mem[4048] = 4'b0000;
	mem[4049] = 4'b0000;
	mem[4050] = 4'b0000;
	mem[4051] = 4'b0000;
	mem[4052] = 4'b0000;
	mem[4053] = 4'b0000;
	mem[4054] = 4'b0000;
	mem[4055] = 4'b0000;
	mem[4056] = 4'b0000;
	mem[4057] = 4'b0000;
	mem[4058] = 4'b0000;
	mem[4059] = 4'b0000;
	mem[4060] = 4'b0000;
	mem[4061] = 4'b0000;
	mem[4062] = 4'b0000;
	mem[4063] = 4'b0000;
	mem[4064] = 4'b0000;
	mem[4065] = 4'b0000;
	mem[4066] = 4'b0000;
	mem[4067] = 4'b0000;
	mem[4068] = 4'b0000;
	mem[4069] = 4'b0000;
	mem[4070] = 4'b0000;
	mem[4071] = 4'b0000;
	mem[4072] = 4'b0000;
	mem[4073] = 4'b0000;
	mem[4074] = 4'b0000;
	mem[4075] = 4'b0000;
	mem[4076] = 4'b0000;
	mem[4077] = 4'b0000;
	mem[4078] = 4'b0000;
	mem[4079] = 4'b0000;
	mem[4080] = 4'b0000;
	mem[4081] = 4'b0000;
	mem[4082] = 4'b0000;
	mem[4083] = 4'b0000;
	mem[4084] = 4'b0000;
	mem[4085] = 4'b0000;
	mem[4086] = 4'b0000;
	mem[4087] = 4'b0000;
	mem[4088] = 4'b0000;
	mem[4089] = 4'b0000;
	mem[4090] = 4'b0000;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_0b (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0000;
	mem[4] = 4'b0000;
	mem[5] = 4'b0000;
	mem[6] = 4'b0000;
	mem[7] = 4'b0000;
	mem[8] = 4'b0000;
	mem[9] = 4'b0000;
	mem[10] = 4'b0000;
	mem[11] = 4'b0000;
	mem[12] = 4'b0000;
	mem[13] = 4'b0000;
	mem[14] = 4'b0000;
	mem[15] = 4'b0000;
	mem[16] = 4'b0000;
	mem[17] = 4'b0000;
	mem[18] = 4'b0000;
	mem[19] = 4'b0000;
	mem[20] = 4'b0000;
	mem[21] = 4'b0000;
	mem[22] = 4'b0000;
	mem[23] = 4'b0000;
	mem[24] = 4'b0000;
	mem[25] = 4'b0000;
	mem[26] = 4'b0000;
	mem[27] = 4'b0000;
	mem[28] = 4'b0000;
	mem[29] = 4'b0000;
	mem[30] = 4'b0000;
	mem[31] = 4'b0000;
	mem[32] = 4'b0000;
	mem[33] = 4'b0000;
	mem[34] = 4'b0000;
	mem[35] = 4'b0000;
	mem[36] = 4'b0000;
	mem[37] = 4'b0000;
	mem[38] = 4'b0000;
	mem[39] = 4'b0000;
	mem[40] = 4'b0000;
	mem[41] = 4'b0000;
	mem[42] = 4'b0000;
	mem[43] = 4'b0000;
	mem[44] = 4'b0000;
	mem[45] = 4'b0000;
	mem[46] = 4'b0000;
	mem[47] = 4'b0000;
	mem[48] = 4'b0000;
	mem[49] = 4'b0000;
	mem[50] = 4'b0000;
	mem[51] = 4'b0000;
	mem[52] = 4'b0000;
	mem[53] = 4'b0000;
	mem[54] = 4'b0000;
	mem[55] = 4'b0000;
	mem[56] = 4'b0000;
	mem[57] = 4'b0000;
	mem[58] = 4'b0000;
	mem[59] = 4'b0000;
	mem[60] = 4'b0000;
	mem[61] = 4'b0000;
	mem[62] = 4'b0000;
	mem[63] = 4'b0000;
	mem[64] = 4'b0000;
	mem[65] = 4'b0000;
	mem[66] = 4'b0000;
	mem[67] = 4'b0000;
	mem[68] = 4'b0000;
	mem[69] = 4'b0000;
	mem[70] = 4'b0000;
	mem[71] = 4'b0000;
	mem[72] = 4'b0000;
	mem[73] = 4'b0000;
	mem[74] = 4'b0000;
	mem[75] = 4'b0000;
	mem[76] = 4'b0000;
	mem[77] = 4'b0000;
	mem[78] = 4'b0000;
	mem[79] = 4'b0000;
	mem[80] = 4'b0000;
	mem[81] = 4'b0000;
	mem[82] = 4'b0000;
	mem[83] = 4'b0000;
	mem[84] = 4'b0000;
	mem[85] = 4'b0000;
	mem[86] = 4'b0000;
	mem[87] = 4'b0000;
	mem[88] = 4'b0000;
	mem[89] = 4'b0000;
	mem[90] = 4'b0000;
	mem[91] = 4'b0000;
	mem[92] = 4'b0000;
	mem[93] = 4'b0000;
	mem[94] = 4'b0000;
	mem[95] = 4'b0000;
	mem[96] = 4'b0000;
	mem[97] = 4'b0000;
	mem[98] = 4'b0000;
	mem[99] = 4'b0000;
	mem[100] = 4'b0000;
	mem[101] = 4'b0000;
	mem[102] = 4'b0000;
	mem[103] = 4'b0000;
	mem[104] = 4'b0000;
	mem[105] = 4'b0000;
	mem[106] = 4'b0000;
	mem[107] = 4'b0000;
	mem[108] = 4'b0000;
	mem[109] = 4'b0000;
	mem[110] = 4'b0000;
	mem[111] = 4'b0000;
	mem[112] = 4'b0000;
	mem[113] = 4'b0000;
	mem[114] = 4'b0000;
	mem[115] = 4'b0000;
	mem[116] = 4'b0000;
	mem[117] = 4'b0000;
	mem[118] = 4'b0000;
	mem[119] = 4'b0000;
	mem[120] = 4'b0000;
	mem[121] = 4'b0000;
	mem[122] = 4'b0000;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b0000;
	mem[132] = 4'b0000;
	mem[133] = 4'b0000;
	mem[134] = 4'b0000;
	mem[135] = 4'b0000;
	mem[136] = 4'b0000;
	mem[137] = 4'b0000;
	mem[138] = 4'b0000;
	mem[139] = 4'b0000;
	mem[140] = 4'b0000;
	mem[141] = 4'b0000;
	mem[142] = 4'b0000;
	mem[143] = 4'b0000;
	mem[144] = 4'b0000;
	mem[145] = 4'b0000;
	mem[146] = 4'b0000;
	mem[147] = 4'b0000;
	mem[148] = 4'b0000;
	mem[149] = 4'b0000;
	mem[150] = 4'b0000;
	mem[151] = 4'b0000;
	mem[152] = 4'b0000;
	mem[153] = 4'b0000;
	mem[154] = 4'b0000;
	mem[155] = 4'b0000;
	mem[156] = 4'b0000;
	mem[157] = 4'b0000;
	mem[158] = 4'b0000;
	mem[159] = 4'b0000;
	mem[160] = 4'b0000;
	mem[161] = 4'b0000;
	mem[162] = 4'b0000;
	mem[163] = 4'b0000;
	mem[164] = 4'b0000;
	mem[165] = 4'b0000;
	mem[166] = 4'b0000;
	mem[167] = 4'b0000;
	mem[168] = 4'b0000;
	mem[169] = 4'b0000;
	mem[170] = 4'b0000;
	mem[171] = 4'b0000;
	mem[172] = 4'b0000;
	mem[173] = 4'b0000;
	mem[174] = 4'b0000;
	mem[175] = 4'b0000;
	mem[176] = 4'b0000;
	mem[177] = 4'b0000;
	mem[178] = 4'b0000;
	mem[179] = 4'b0000;
	mem[180] = 4'b0000;
	mem[181] = 4'b0000;
	mem[182] = 4'b0000;
	mem[183] = 4'b0000;
	mem[184] = 4'b0000;
	mem[185] = 4'b0000;
	mem[186] = 4'b0000;
	mem[187] = 4'b0000;
	mem[188] = 4'b0000;
	mem[189] = 4'b0000;
	mem[190] = 4'b0000;
	mem[191] = 4'b0000;
	mem[192] = 4'b0000;
	mem[193] = 4'b0000;
	mem[194] = 4'b0000;
	mem[195] = 4'b0000;
	mem[196] = 4'b0000;
	mem[197] = 4'b0000;
	mem[198] = 4'b0000;
	mem[199] = 4'b0000;
	mem[200] = 4'b0000;
	mem[201] = 4'b0000;
	mem[202] = 4'b0000;
	mem[203] = 4'b0000;
	mem[204] = 4'b0000;
	mem[205] = 4'b0000;
	mem[206] = 4'b0000;
	mem[207] = 4'b0000;
	mem[208] = 4'b0000;
	mem[209] = 4'b0000;
	mem[210] = 4'b0000;
	mem[211] = 4'b0000;
	mem[212] = 4'b0000;
	mem[213] = 4'b0000;
	mem[214] = 4'b0000;
	mem[215] = 4'b0000;
	mem[216] = 4'b0000;
	mem[217] = 4'b0000;
	mem[218] = 4'b0000;
	mem[219] = 4'b0000;
	mem[220] = 4'b0000;
	mem[221] = 4'b0000;
	mem[222] = 4'b0000;
	mem[223] = 4'b0000;
	mem[224] = 4'b0000;
	mem[225] = 4'b0000;
	mem[226] = 4'b0000;
	mem[227] = 4'b0000;
	mem[228] = 4'b0000;
	mem[229] = 4'b0000;
	mem[230] = 4'b0000;
	mem[231] = 4'b0000;
	mem[232] = 4'b0000;
	mem[233] = 4'b0000;
	mem[234] = 4'b0000;
	mem[235] = 4'b0000;
	mem[236] = 4'b0000;
	mem[237] = 4'b0000;
	mem[238] = 4'b0000;
	mem[239] = 4'b0000;
	mem[240] = 4'b0000;
	mem[241] = 4'b0000;
	mem[242] = 4'b0000;
	mem[243] = 4'b0000;
	mem[244] = 4'b0000;
	mem[245] = 4'b0000;
	mem[246] = 4'b0000;
	mem[247] = 4'b0000;
	mem[248] = 4'b0000;
	mem[249] = 4'b0000;
	mem[250] = 4'b0000;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0000;
	mem[260] = 4'b0000;
	mem[261] = 4'b0000;
	mem[262] = 4'b0000;
	mem[263] = 4'b0000;
	mem[264] = 4'b0000;
	mem[265] = 4'b0000;
	mem[266] = 4'b0000;
	mem[267] = 4'b0000;
	mem[268] = 4'b0000;
	mem[269] = 4'b0000;
	mem[270] = 4'b0000;
	mem[271] = 4'b0000;
	mem[272] = 4'b0000;
	mem[273] = 4'b0000;
	mem[274] = 4'b0000;
	mem[275] = 4'b0000;
	mem[276] = 4'b0000;
	mem[277] = 4'b0000;
	mem[278] = 4'b0000;
	mem[279] = 4'b0000;
	mem[280] = 4'b0000;
	mem[281] = 4'b0000;
	mem[282] = 4'b0000;
	mem[283] = 4'b0000;
	mem[284] = 4'b0000;
	mem[285] = 4'b0000;
	mem[286] = 4'b0000;
	mem[287] = 4'b0000;
	mem[288] = 4'b0000;
	mem[289] = 4'b0000;
	mem[290] = 4'b0000;
	mem[291] = 4'b0000;
	mem[292] = 4'b0000;
	mem[293] = 4'b0000;
	mem[294] = 4'b0000;
	mem[295] = 4'b0000;
	mem[296] = 4'b0000;
	mem[297] = 4'b0000;
	mem[298] = 4'b0000;
	mem[299] = 4'b0000;
	mem[300] = 4'b0000;
	mem[301] = 4'b0000;
	mem[302] = 4'b0000;
	mem[303] = 4'b0000;
	mem[304] = 4'b0000;
	mem[305] = 4'b0000;
	mem[306] = 4'b0000;
	mem[307] = 4'b0000;
	mem[308] = 4'b0000;
	mem[309] = 4'b0000;
	mem[310] = 4'b0000;
	mem[311] = 4'b0000;
	mem[312] = 4'b0000;
	mem[313] = 4'b0000;
	mem[314] = 4'b0000;
	mem[315] = 4'b0000;
	mem[316] = 4'b0000;
	mem[317] = 4'b0000;
	mem[318] = 4'b0000;
	mem[319] = 4'b0000;
	mem[320] = 4'b0000;
	mem[321] = 4'b0000;
	mem[322] = 4'b0000;
	mem[323] = 4'b0000;
	mem[324] = 4'b0000;
	mem[325] = 4'b0000;
	mem[326] = 4'b0000;
	mem[327] = 4'b0000;
	mem[328] = 4'b0000;
	mem[329] = 4'b0000;
	mem[330] = 4'b0000;
	mem[331] = 4'b0000;
	mem[332] = 4'b0000;
	mem[333] = 4'b0000;
	mem[334] = 4'b0000;
	mem[335] = 4'b0000;
	mem[336] = 4'b0000;
	mem[337] = 4'b0000;
	mem[338] = 4'b0000;
	mem[339] = 4'b0000;
	mem[340] = 4'b0000;
	mem[341] = 4'b0000;
	mem[342] = 4'b0000;
	mem[343] = 4'b0000;
	mem[344] = 4'b0000;
	mem[345] = 4'b0000;
	mem[346] = 4'b0000;
	mem[347] = 4'b0000;
	mem[348] = 4'b0000;
	mem[349] = 4'b0000;
	mem[350] = 4'b0000;
	mem[351] = 4'b0000;
	mem[352] = 4'b0000;
	mem[353] = 4'b0000;
	mem[354] = 4'b0000;
	mem[355] = 4'b0000;
	mem[356] = 4'b0000;
	mem[357] = 4'b0000;
	mem[358] = 4'b0000;
	mem[359] = 4'b0000;
	mem[360] = 4'b0000;
	mem[361] = 4'b0000;
	mem[362] = 4'b0000;
	mem[363] = 4'b0000;
	mem[364] = 4'b0000;
	mem[365] = 4'b0000;
	mem[366] = 4'b0000;
	mem[367] = 4'b0000;
	mem[368] = 4'b0000;
	mem[369] = 4'b0000;
	mem[370] = 4'b0000;
	mem[371] = 4'b0000;
	mem[372] = 4'b0000;
	mem[373] = 4'b0000;
	mem[374] = 4'b0000;
	mem[375] = 4'b0000;
	mem[376] = 4'b0000;
	mem[377] = 4'b0000;
	mem[378] = 4'b0000;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0000;
	mem[388] = 4'b0000;
	mem[389] = 4'b0000;
	mem[390] = 4'b0000;
	mem[391] = 4'b0000;
	mem[392] = 4'b0000;
	mem[393] = 4'b0000;
	mem[394] = 4'b0000;
	mem[395] = 4'b0000;
	mem[396] = 4'b0000;
	mem[397] = 4'b0000;
	mem[398] = 4'b0000;
	mem[399] = 4'b0000;
	mem[400] = 4'b0000;
	mem[401] = 4'b0000;
	mem[402] = 4'b0000;
	mem[403] = 4'b0000;
	mem[404] = 4'b0000;
	mem[405] = 4'b0000;
	mem[406] = 4'b0000;
	mem[407] = 4'b0000;
	mem[408] = 4'b0000;
	mem[409] = 4'b0000;
	mem[410] = 4'b0000;
	mem[411] = 4'b0000;
	mem[412] = 4'b0000;
	mem[413] = 4'b0000;
	mem[414] = 4'b0000;
	mem[415] = 4'b0000;
	mem[416] = 4'b0000;
	mem[417] = 4'b0000;
	mem[418] = 4'b0000;
	mem[419] = 4'b0000;
	mem[420] = 4'b0000;
	mem[421] = 4'b0000;
	mem[422] = 4'b0000;
	mem[423] = 4'b0000;
	mem[424] = 4'b0000;
	mem[425] = 4'b0000;
	mem[426] = 4'b0000;
	mem[427] = 4'b0000;
	mem[428] = 4'b0000;
	mem[429] = 4'b0000;
	mem[430] = 4'b0000;
	mem[431] = 4'b0000;
	mem[432] = 4'b0000;
	mem[433] = 4'b0000;
	mem[434] = 4'b0000;
	mem[435] = 4'b0000;
	mem[436] = 4'b0000;
	mem[437] = 4'b0000;
	mem[438] = 4'b0000;
	mem[439] = 4'b0000;
	mem[440] = 4'b0000;
	mem[441] = 4'b0000;
	mem[442] = 4'b0000;
	mem[443] = 4'b0000;
	mem[444] = 4'b0000;
	mem[445] = 4'b0000;
	mem[446] = 4'b0000;
	mem[447] = 4'b0000;
	mem[448] = 4'b0000;
	mem[449] = 4'b0000;
	mem[450] = 4'b0000;
	mem[451] = 4'b0000;
	mem[452] = 4'b0000;
	mem[453] = 4'b0000;
	mem[454] = 4'b0000;
	mem[455] = 4'b0000;
	mem[456] = 4'b0000;
	mem[457] = 4'b0000;
	mem[458] = 4'b0000;
	mem[459] = 4'b0000;
	mem[460] = 4'b0000;
	mem[461] = 4'b0000;
	mem[462] = 4'b0000;
	mem[463] = 4'b0000;
	mem[464] = 4'b0000;
	mem[465] = 4'b0000;
	mem[466] = 4'b0000;
	mem[467] = 4'b0000;
	mem[468] = 4'b0000;
	mem[469] = 4'b0000;
	mem[470] = 4'b0000;
	mem[471] = 4'b0000;
	mem[472] = 4'b0000;
	mem[473] = 4'b0000;
	mem[474] = 4'b0000;
	mem[475] = 4'b0000;
	mem[476] = 4'b0000;
	mem[477] = 4'b0000;
	mem[478] = 4'b0000;
	mem[479] = 4'b0000;
	mem[480] = 4'b0000;
	mem[481] = 4'b0000;
	mem[482] = 4'b0000;
	mem[483] = 4'b0000;
	mem[484] = 4'b0000;
	mem[485] = 4'b0000;
	mem[486] = 4'b0000;
	mem[487] = 4'b0000;
	mem[488] = 4'b0000;
	mem[489] = 4'b0000;
	mem[490] = 4'b0000;
	mem[491] = 4'b0000;
	mem[492] = 4'b0000;
	mem[493] = 4'b0000;
	mem[494] = 4'b0000;
	mem[495] = 4'b0000;
	mem[496] = 4'b0000;
	mem[497] = 4'b0000;
	mem[498] = 4'b0000;
	mem[499] = 4'b0000;
	mem[500] = 4'b0000;
	mem[501] = 4'b0000;
	mem[502] = 4'b0000;
	mem[503] = 4'b0000;
	mem[504] = 4'b0000;
	mem[505] = 4'b0000;
	mem[506] = 4'b0000;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0000;
	mem[516] = 4'b0000;
	mem[517] = 4'b0000;
	mem[518] = 4'b0000;
	mem[519] = 4'b0000;
	mem[520] = 4'b0000;
	mem[521] = 4'b0000;
	mem[522] = 4'b0000;
	mem[523] = 4'b0000;
	mem[524] = 4'b0000;
	mem[525] = 4'b0000;
	mem[526] = 4'b0000;
	mem[527] = 4'b0000;
	mem[528] = 4'b0000;
	mem[529] = 4'b0000;
	mem[530] = 4'b0000;
	mem[531] = 4'b0000;
	mem[532] = 4'b0000;
	mem[533] = 4'b0000;
	mem[534] = 4'b0000;
	mem[535] = 4'b0000;
	mem[536] = 4'b0000;
	mem[537] = 4'b0000;
	mem[538] = 4'b0000;
	mem[539] = 4'b0000;
	mem[540] = 4'b0000;
	mem[541] = 4'b0000;
	mem[542] = 4'b0000;
	mem[543] = 4'b0000;
	mem[544] = 4'b0000;
	mem[545] = 4'b0000;
	mem[546] = 4'b0000;
	mem[547] = 4'b0000;
	mem[548] = 4'b0000;
	mem[549] = 4'b0000;
	mem[550] = 4'b0000;
	mem[551] = 4'b0000;
	mem[552] = 4'b0000;
	mem[553] = 4'b0000;
	mem[554] = 4'b0000;
	mem[555] = 4'b0000;
	mem[556] = 4'b0000;
	mem[557] = 4'b0000;
	mem[558] = 4'b0000;
	mem[559] = 4'b0000;
	mem[560] = 4'b0000;
	mem[561] = 4'b0000;
	mem[562] = 4'b0000;
	mem[563] = 4'b0000;
	mem[564] = 4'b0000;
	mem[565] = 4'b0000;
	mem[566] = 4'b0000;
	mem[567] = 4'b0000;
	mem[568] = 4'b0000;
	mem[569] = 4'b0000;
	mem[570] = 4'b0000;
	mem[571] = 4'b0000;
	mem[572] = 4'b0000;
	mem[573] = 4'b0000;
	mem[574] = 4'b0000;
	mem[575] = 4'b0000;
	mem[576] = 4'b0000;
	mem[577] = 4'b0000;
	mem[578] = 4'b0000;
	mem[579] = 4'b0000;
	mem[580] = 4'b0000;
	mem[581] = 4'b0000;
	mem[582] = 4'b0000;
	mem[583] = 4'b0000;
	mem[584] = 4'b0000;
	mem[585] = 4'b0000;
	mem[586] = 4'b0000;
	mem[587] = 4'b0000;
	mem[588] = 4'b0000;
	mem[589] = 4'b0000;
	mem[590] = 4'b0000;
	mem[591] = 4'b0000;
	mem[592] = 4'b0000;
	mem[593] = 4'b0000;
	mem[594] = 4'b0000;
	mem[595] = 4'b0000;
	mem[596] = 4'b0000;
	mem[597] = 4'b0000;
	mem[598] = 4'b0000;
	mem[599] = 4'b0000;
	mem[600] = 4'b0000;
	mem[601] = 4'b0000;
	mem[602] = 4'b0000;
	mem[603] = 4'b0000;
	mem[604] = 4'b0000;
	mem[605] = 4'b0000;
	mem[606] = 4'b0000;
	mem[607] = 4'b0000;
	mem[608] = 4'b0000;
	mem[609] = 4'b0000;
	mem[610] = 4'b0000;
	mem[611] = 4'b0000;
	mem[612] = 4'b0000;
	mem[613] = 4'b0000;
	mem[614] = 4'b0000;
	mem[615] = 4'b0000;
	mem[616] = 4'b0000;
	mem[617] = 4'b0000;
	mem[618] = 4'b0000;
	mem[619] = 4'b0000;
	mem[620] = 4'b0000;
	mem[621] = 4'b0000;
	mem[622] = 4'b0000;
	mem[623] = 4'b0000;
	mem[624] = 4'b0000;
	mem[625] = 4'b0000;
	mem[626] = 4'b0000;
	mem[627] = 4'b0000;
	mem[628] = 4'b0000;
	mem[629] = 4'b0000;
	mem[630] = 4'b0000;
	mem[631] = 4'b0000;
	mem[632] = 4'b0000;
	mem[633] = 4'b0000;
	mem[634] = 4'b0000;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0000;
	mem[644] = 4'b0000;
	mem[645] = 4'b0000;
	mem[646] = 4'b0000;
	mem[647] = 4'b0000;
	mem[648] = 4'b0000;
	mem[649] = 4'b0000;
	mem[650] = 4'b0000;
	mem[651] = 4'b0000;
	mem[652] = 4'b0000;
	mem[653] = 4'b0000;
	mem[654] = 4'b0000;
	mem[655] = 4'b0000;
	mem[656] = 4'b0000;
	mem[657] = 4'b0000;
	mem[658] = 4'b0000;
	mem[659] = 4'b0000;
	mem[660] = 4'b0000;
	mem[661] = 4'b0000;
	mem[662] = 4'b0000;
	mem[663] = 4'b0000;
	mem[664] = 4'b0000;
	mem[665] = 4'b0000;
	mem[666] = 4'b0000;
	mem[667] = 4'b0000;
	mem[668] = 4'b0000;
	mem[669] = 4'b0000;
	mem[670] = 4'b0000;
	mem[671] = 4'b0000;
	mem[672] = 4'b0000;
	mem[673] = 4'b0000;
	mem[674] = 4'b0000;
	mem[675] = 4'b0000;
	mem[676] = 4'b0000;
	mem[677] = 4'b0000;
	mem[678] = 4'b0000;
	mem[679] = 4'b0000;
	mem[680] = 4'b0000;
	mem[681] = 4'b0000;
	mem[682] = 4'b0000;
	mem[683] = 4'b0000;
	mem[684] = 4'b0000;
	mem[685] = 4'b0000;
	mem[686] = 4'b0000;
	mem[687] = 4'b0000;
	mem[688] = 4'b0000;
	mem[689] = 4'b0000;
	mem[690] = 4'b0000;
	mem[691] = 4'b0000;
	mem[692] = 4'b0000;
	mem[693] = 4'b0000;
	mem[694] = 4'b0000;
	mem[695] = 4'b0000;
	mem[696] = 4'b0000;
	mem[697] = 4'b0000;
	mem[698] = 4'b0000;
	mem[699] = 4'b0000;
	mem[700] = 4'b0000;
	mem[701] = 4'b0000;
	mem[702] = 4'b0000;
	mem[703] = 4'b0000;
	mem[704] = 4'b0000;
	mem[705] = 4'b0000;
	mem[706] = 4'b0000;
	mem[707] = 4'b0000;
	mem[708] = 4'b0000;
	mem[709] = 4'b0000;
	mem[710] = 4'b0000;
	mem[711] = 4'b0000;
	mem[712] = 4'b0000;
	mem[713] = 4'b0000;
	mem[714] = 4'b0000;
	mem[715] = 4'b0000;
	mem[716] = 4'b0000;
	mem[717] = 4'b0000;
	mem[718] = 4'b0000;
	mem[719] = 4'b0000;
	mem[720] = 4'b0000;
	mem[721] = 4'b0000;
	mem[722] = 4'b0000;
	mem[723] = 4'b0000;
	mem[724] = 4'b0000;
	mem[725] = 4'b0000;
	mem[726] = 4'b0000;
	mem[727] = 4'b0000;
	mem[728] = 4'b0000;
	mem[729] = 4'b0000;
	mem[730] = 4'b0000;
	mem[731] = 4'b0000;
	mem[732] = 4'b0000;
	mem[733] = 4'b0000;
	mem[734] = 4'b0000;
	mem[735] = 4'b0000;
	mem[736] = 4'b0000;
	mem[737] = 4'b0000;
	mem[738] = 4'b0000;
	mem[739] = 4'b0000;
	mem[740] = 4'b0000;
	mem[741] = 4'b0000;
	mem[742] = 4'b0000;
	mem[743] = 4'b0000;
	mem[744] = 4'b0000;
	mem[745] = 4'b0000;
	mem[746] = 4'b0000;
	mem[747] = 4'b0000;
	mem[748] = 4'b0000;
	mem[749] = 4'b0000;
	mem[750] = 4'b0000;
	mem[751] = 4'b0000;
	mem[752] = 4'b0000;
	mem[753] = 4'b0000;
	mem[754] = 4'b0000;
	mem[755] = 4'b0000;
	mem[756] = 4'b0000;
	mem[757] = 4'b0000;
	mem[758] = 4'b0000;
	mem[759] = 4'b0000;
	mem[760] = 4'b0000;
	mem[761] = 4'b0000;
	mem[762] = 4'b0000;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0000;
	mem[772] = 4'b0000;
	mem[773] = 4'b0000;
	mem[774] = 4'b0000;
	mem[775] = 4'b0000;
	mem[776] = 4'b0000;
	mem[777] = 4'b0000;
	mem[778] = 4'b0000;
	mem[779] = 4'b0000;
	mem[780] = 4'b0000;
	mem[781] = 4'b0000;
	mem[782] = 4'b0000;
	mem[783] = 4'b0000;
	mem[784] = 4'b0000;
	mem[785] = 4'b0000;
	mem[786] = 4'b0000;
	mem[787] = 4'b0000;
	mem[788] = 4'b0000;
	mem[789] = 4'b0000;
	mem[790] = 4'b0000;
	mem[791] = 4'b0000;
	mem[792] = 4'b0000;
	mem[793] = 4'b0000;
	mem[794] = 4'b0000;
	mem[795] = 4'b0000;
	mem[796] = 4'b0000;
	mem[797] = 4'b0000;
	mem[798] = 4'b0000;
	mem[799] = 4'b0000;
	mem[800] = 4'b0000;
	mem[801] = 4'b0000;
	mem[802] = 4'b0000;
	mem[803] = 4'b0000;
	mem[804] = 4'b0000;
	mem[805] = 4'b0000;
	mem[806] = 4'b0000;
	mem[807] = 4'b0000;
	mem[808] = 4'b0000;
	mem[809] = 4'b0000;
	mem[810] = 4'b0000;
	mem[811] = 4'b0000;
	mem[812] = 4'b0000;
	mem[813] = 4'b0000;
	mem[814] = 4'b0000;
	mem[815] = 4'b0000;
	mem[816] = 4'b0000;
	mem[817] = 4'b0000;
	mem[818] = 4'b0000;
	mem[819] = 4'b0000;
	mem[820] = 4'b0000;
	mem[821] = 4'b0000;
	mem[822] = 4'b0000;
	mem[823] = 4'b0000;
	mem[824] = 4'b0000;
	mem[825] = 4'b0000;
	mem[826] = 4'b0000;
	mem[827] = 4'b0000;
	mem[828] = 4'b0000;
	mem[829] = 4'b0000;
	mem[830] = 4'b0000;
	mem[831] = 4'b0000;
	mem[832] = 4'b0000;
	mem[833] = 4'b0000;
	mem[834] = 4'b0000;
	mem[835] = 4'b0000;
	mem[836] = 4'b0000;
	mem[837] = 4'b0000;
	mem[838] = 4'b0000;
	mem[839] = 4'b0000;
	mem[840] = 4'b0000;
	mem[841] = 4'b0000;
	mem[842] = 4'b0000;
	mem[843] = 4'b0000;
	mem[844] = 4'b0000;
	mem[845] = 4'b0000;
	mem[846] = 4'b0000;
	mem[847] = 4'b0000;
	mem[848] = 4'b0000;
	mem[849] = 4'b0000;
	mem[850] = 4'b0000;
	mem[851] = 4'b0000;
	mem[852] = 4'b0000;
	mem[853] = 4'b0000;
	mem[854] = 4'b0000;
	mem[855] = 4'b0000;
	mem[856] = 4'b0000;
	mem[857] = 4'b0000;
	mem[858] = 4'b0000;
	mem[859] = 4'b0000;
	mem[860] = 4'b0000;
	mem[861] = 4'b0000;
	mem[862] = 4'b0000;
	mem[863] = 4'b0000;
	mem[864] = 4'b0000;
	mem[865] = 4'b0000;
	mem[866] = 4'b0000;
	mem[867] = 4'b0000;
	mem[868] = 4'b0000;
	mem[869] = 4'b0000;
	mem[870] = 4'b0000;
	mem[871] = 4'b0000;
	mem[872] = 4'b0000;
	mem[873] = 4'b0000;
	mem[874] = 4'b0000;
	mem[875] = 4'b0000;
	mem[876] = 4'b0000;
	mem[877] = 4'b0000;
	mem[878] = 4'b0000;
	mem[879] = 4'b0000;
	mem[880] = 4'b0000;
	mem[881] = 4'b0000;
	mem[882] = 4'b0000;
	mem[883] = 4'b0000;
	mem[884] = 4'b0000;
	mem[885] = 4'b0000;
	mem[886] = 4'b0000;
	mem[887] = 4'b0000;
	mem[888] = 4'b0000;
	mem[889] = 4'b0000;
	mem[890] = 4'b0000;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0000;
	mem[900] = 4'b0000;
	mem[901] = 4'b0000;
	mem[902] = 4'b0000;
	mem[903] = 4'b0000;
	mem[904] = 4'b0000;
	mem[905] = 4'b0000;
	mem[906] = 4'b0000;
	mem[907] = 4'b0000;
	mem[908] = 4'b0000;
	mem[909] = 4'b0000;
	mem[910] = 4'b0000;
	mem[911] = 4'b0000;
	mem[912] = 4'b0000;
	mem[913] = 4'b0000;
	mem[914] = 4'b0000;
	mem[915] = 4'b0000;
	mem[916] = 4'b0000;
	mem[917] = 4'b0000;
	mem[918] = 4'b0000;
	mem[919] = 4'b0000;
	mem[920] = 4'b0000;
	mem[921] = 4'b0000;
	mem[922] = 4'b0000;
	mem[923] = 4'b0000;
	mem[924] = 4'b0000;
	mem[925] = 4'b0000;
	mem[926] = 4'b0000;
	mem[927] = 4'b0000;
	mem[928] = 4'b0000;
	mem[929] = 4'b0000;
	mem[930] = 4'b0000;
	mem[931] = 4'b0000;
	mem[932] = 4'b0000;
	mem[933] = 4'b0000;
	mem[934] = 4'b0000;
	mem[935] = 4'b0000;
	mem[936] = 4'b0000;
	mem[937] = 4'b0000;
	mem[938] = 4'b0000;
	mem[939] = 4'b0000;
	mem[940] = 4'b0000;
	mem[941] = 4'b0000;
	mem[942] = 4'b0000;
	mem[943] = 4'b0000;
	mem[944] = 4'b0000;
	mem[945] = 4'b0000;
	mem[946] = 4'b0000;
	mem[947] = 4'b0000;
	mem[948] = 4'b0000;
	mem[949] = 4'b0000;
	mem[950] = 4'b0000;
	mem[951] = 4'b0000;
	mem[952] = 4'b0000;
	mem[953] = 4'b0000;
	mem[954] = 4'b0000;
	mem[955] = 4'b0000;
	mem[956] = 4'b0000;
	mem[957] = 4'b0000;
	mem[958] = 4'b0000;
	mem[959] = 4'b0000;
	mem[960] = 4'b0000;
	mem[961] = 4'b0000;
	mem[962] = 4'b0000;
	mem[963] = 4'b0000;
	mem[964] = 4'b0000;
	mem[965] = 4'b0000;
	mem[966] = 4'b0000;
	mem[967] = 4'b0000;
	mem[968] = 4'b0000;
	mem[969] = 4'b0000;
	mem[970] = 4'b0000;
	mem[971] = 4'b0000;
	mem[972] = 4'b0000;
	mem[973] = 4'b0000;
	mem[974] = 4'b0000;
	mem[975] = 4'b0000;
	mem[976] = 4'b0000;
	mem[977] = 4'b0000;
	mem[978] = 4'b0000;
	mem[979] = 4'b0000;
	mem[980] = 4'b0000;
	mem[981] = 4'b0000;
	mem[982] = 4'b0000;
	mem[983] = 4'b0000;
	mem[984] = 4'b0000;
	mem[985] = 4'b0000;
	mem[986] = 4'b0000;
	mem[987] = 4'b0000;
	mem[988] = 4'b0000;
	mem[989] = 4'b0000;
	mem[990] = 4'b0000;
	mem[991] = 4'b0000;
	mem[992] = 4'b0000;
	mem[993] = 4'b0000;
	mem[994] = 4'b0000;
	mem[995] = 4'b0000;
	mem[996] = 4'b0000;
	mem[997] = 4'b0000;
	mem[998] = 4'b0000;
	mem[999] = 4'b0000;
	mem[1000] = 4'b0000;
	mem[1001] = 4'b0000;
	mem[1002] = 4'b0000;
	mem[1003] = 4'b0000;
	mem[1004] = 4'b0000;
	mem[1005] = 4'b0000;
	mem[1006] = 4'b0000;
	mem[1007] = 4'b0000;
	mem[1008] = 4'b0000;
	mem[1009] = 4'b0000;
	mem[1010] = 4'b0000;
	mem[1011] = 4'b0000;
	mem[1012] = 4'b0000;
	mem[1013] = 4'b0000;
	mem[1014] = 4'b0000;
	mem[1015] = 4'b0000;
	mem[1016] = 4'b0000;
	mem[1017] = 4'b0000;
	mem[1018] = 4'b0000;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0000;
	mem[1028] = 4'b0000;
	mem[1029] = 4'b0000;
	mem[1030] = 4'b0000;
	mem[1031] = 4'b0000;
	mem[1032] = 4'b0000;
	mem[1033] = 4'b0000;
	mem[1034] = 4'b0000;
	mem[1035] = 4'b0000;
	mem[1036] = 4'b0000;
	mem[1037] = 4'b0000;
	mem[1038] = 4'b0000;
	mem[1039] = 4'b0000;
	mem[1040] = 4'b0000;
	mem[1041] = 4'b0000;
	mem[1042] = 4'b0000;
	mem[1043] = 4'b0000;
	mem[1044] = 4'b0000;
	mem[1045] = 4'b0000;
	mem[1046] = 4'b0000;
	mem[1047] = 4'b0000;
	mem[1048] = 4'b0000;
	mem[1049] = 4'b0000;
	mem[1050] = 4'b0000;
	mem[1051] = 4'b0000;
	mem[1052] = 4'b0000;
	mem[1053] = 4'b0000;
	mem[1054] = 4'b0000;
	mem[1055] = 4'b0000;
	mem[1056] = 4'b0000;
	mem[1057] = 4'b0000;
	mem[1058] = 4'b0000;
	mem[1059] = 4'b0000;
	mem[1060] = 4'b0000;
	mem[1061] = 4'b0000;
	mem[1062] = 4'b0000;
	mem[1063] = 4'b0000;
	mem[1064] = 4'b0000;
	mem[1065] = 4'b0000;
	mem[1066] = 4'b0000;
	mem[1067] = 4'b0000;
	mem[1068] = 4'b0000;
	mem[1069] = 4'b0000;
	mem[1070] = 4'b0000;
	mem[1071] = 4'b0000;
	mem[1072] = 4'b0000;
	mem[1073] = 4'b0000;
	mem[1074] = 4'b0000;
	mem[1075] = 4'b0000;
	mem[1076] = 4'b0000;
	mem[1077] = 4'b0000;
	mem[1078] = 4'b0000;
	mem[1079] = 4'b0000;
	mem[1080] = 4'b0000;
	mem[1081] = 4'b0000;
	mem[1082] = 4'b0000;
	mem[1083] = 4'b0000;
	mem[1084] = 4'b0000;
	mem[1085] = 4'b0000;
	mem[1086] = 4'b0000;
	mem[1087] = 4'b0000;
	mem[1088] = 4'b0000;
	mem[1089] = 4'b0001;
	mem[1090] = 4'b0001;
	mem[1091] = 4'b0000;
	mem[1092] = 4'b0000;
	mem[1093] = 4'b0000;
	mem[1094] = 4'b0000;
	mem[1095] = 4'b0000;
	mem[1096] = 4'b0000;
	mem[1097] = 4'b0000;
	mem[1098] = 4'b0000;
	mem[1099] = 4'b0000;
	mem[1100] = 4'b0000;
	mem[1101] = 4'b0000;
	mem[1102] = 4'b0000;
	mem[1103] = 4'b0000;
	mem[1104] = 4'b0000;
	mem[1105] = 4'b0000;
	mem[1106] = 4'b0000;
	mem[1107] = 4'b0000;
	mem[1108] = 4'b0000;
	mem[1109] = 4'b0000;
	mem[1110] = 4'b0000;
	mem[1111] = 4'b0000;
	mem[1112] = 4'b0000;
	mem[1113] = 4'b0000;
	mem[1114] = 4'b0000;
	mem[1115] = 4'b0000;
	mem[1116] = 4'b0000;
	mem[1117] = 4'b0000;
	mem[1118] = 4'b0000;
	mem[1119] = 4'b0000;
	mem[1120] = 4'b0000;
	mem[1121] = 4'b0000;
	mem[1122] = 4'b0000;
	mem[1123] = 4'b0000;
	mem[1124] = 4'b0000;
	mem[1125] = 4'b0000;
	mem[1126] = 4'b0000;
	mem[1127] = 4'b0000;
	mem[1128] = 4'b0000;
	mem[1129] = 4'b0000;
	mem[1130] = 4'b0000;
	mem[1131] = 4'b0000;
	mem[1132] = 4'b0000;
	mem[1133] = 4'b0000;
	mem[1134] = 4'b0000;
	mem[1135] = 4'b0000;
	mem[1136] = 4'b0000;
	mem[1137] = 4'b0000;
	mem[1138] = 4'b0000;
	mem[1139] = 4'b0000;
	mem[1140] = 4'b0000;
	mem[1141] = 4'b0000;
	mem[1142] = 4'b0000;
	mem[1143] = 4'b0000;
	mem[1144] = 4'b0000;
	mem[1145] = 4'b0000;
	mem[1146] = 4'b0000;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0000;
	mem[1156] = 4'b0000;
	mem[1157] = 4'b0000;
	mem[1158] = 4'b0000;
	mem[1159] = 4'b0000;
	mem[1160] = 4'b0000;
	mem[1161] = 4'b0000;
	mem[1162] = 4'b0000;
	mem[1163] = 4'b0000;
	mem[1164] = 4'b0000;
	mem[1165] = 4'b0000;
	mem[1166] = 4'b0000;
	mem[1167] = 4'b0000;
	mem[1168] = 4'b0000;
	mem[1169] = 4'b0000;
	mem[1170] = 4'b0000;
	mem[1171] = 4'b0000;
	mem[1172] = 4'b0000;
	mem[1173] = 4'b0000;
	mem[1174] = 4'b0000;
	mem[1175] = 4'b0000;
	mem[1176] = 4'b0000;
	mem[1177] = 4'b0000;
	mem[1178] = 4'b0000;
	mem[1179] = 4'b0000;
	mem[1180] = 4'b0000;
	mem[1181] = 4'b0000;
	mem[1182] = 4'b0000;
	mem[1183] = 4'b0000;
	mem[1184] = 4'b0000;
	mem[1185] = 4'b0000;
	mem[1186] = 4'b0000;
	mem[1187] = 4'b0000;
	mem[1188] = 4'b0000;
	mem[1189] = 4'b0000;
	mem[1190] = 4'b0000;
	mem[1191] = 4'b0000;
	mem[1192] = 4'b0000;
	mem[1193] = 4'b0000;
	mem[1194] = 4'b0000;
	mem[1195] = 4'b0000;
	mem[1196] = 4'b0000;
	mem[1197] = 4'b0000;
	mem[1198] = 4'b0000;
	mem[1199] = 4'b0000;
	mem[1200] = 4'b0000;
	mem[1201] = 4'b0000;
	mem[1202] = 4'b0000;
	mem[1203] = 4'b0000;
	mem[1204] = 4'b0000;
	mem[1205] = 4'b0000;
	mem[1206] = 4'b0000;
	mem[1207] = 4'b0000;
	mem[1208] = 4'b0000;
	mem[1209] = 4'b0000;
	mem[1210] = 4'b0000;
	mem[1211] = 4'b0000;
	mem[1212] = 4'b0000;
	mem[1213] = 4'b0000;
	mem[1214] = 4'b0000;
	mem[1215] = 4'b0000;
	mem[1216] = 4'b0001;
	mem[1217] = 4'b0001;
	mem[1218] = 4'b0000;
	mem[1219] = 4'b0000;
	mem[1220] = 4'b0000;
	mem[1221] = 4'b0000;
	mem[1222] = 4'b0000;
	mem[1223] = 4'b0000;
	mem[1224] = 4'b0000;
	mem[1225] = 4'b0000;
	mem[1226] = 4'b0000;
	mem[1227] = 4'b0000;
	mem[1228] = 4'b0000;
	mem[1229] = 4'b0000;
	mem[1230] = 4'b0000;
	mem[1231] = 4'b0000;
	mem[1232] = 4'b0000;
	mem[1233] = 4'b0000;
	mem[1234] = 4'b0000;
	mem[1235] = 4'b0000;
	mem[1236] = 4'b0000;
	mem[1237] = 4'b0000;
	mem[1238] = 4'b0000;
	mem[1239] = 4'b0000;
	mem[1240] = 4'b0000;
	mem[1241] = 4'b0000;
	mem[1242] = 4'b0000;
	mem[1243] = 4'b0000;
	mem[1244] = 4'b0000;
	mem[1245] = 4'b0000;
	mem[1246] = 4'b0000;
	mem[1247] = 4'b0000;
	mem[1248] = 4'b0000;
	mem[1249] = 4'b0000;
	mem[1250] = 4'b0000;
	mem[1251] = 4'b0000;
	mem[1252] = 4'b0000;
	mem[1253] = 4'b0000;
	mem[1254] = 4'b0000;
	mem[1255] = 4'b0000;
	mem[1256] = 4'b0000;
	mem[1257] = 4'b0000;
	mem[1258] = 4'b0000;
	mem[1259] = 4'b0000;
	mem[1260] = 4'b0000;
	mem[1261] = 4'b0000;
	mem[1262] = 4'b0000;
	mem[1263] = 4'b0000;
	mem[1264] = 4'b0000;
	mem[1265] = 4'b0000;
	mem[1266] = 4'b0000;
	mem[1267] = 4'b0000;
	mem[1268] = 4'b0000;
	mem[1269] = 4'b0000;
	mem[1270] = 4'b0000;
	mem[1271] = 4'b0000;
	mem[1272] = 4'b0000;
	mem[1273] = 4'b0000;
	mem[1274] = 4'b0000;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0000;
	mem[1284] = 4'b0000;
	mem[1285] = 4'b0000;
	mem[1286] = 4'b0000;
	mem[1287] = 4'b0000;
	mem[1288] = 4'b0000;
	mem[1289] = 4'b0000;
	mem[1290] = 4'b0000;
	mem[1291] = 4'b0000;
	mem[1292] = 4'b0000;
	mem[1293] = 4'b0000;
	mem[1294] = 4'b0000;
	mem[1295] = 4'b0000;
	mem[1296] = 4'b0000;
	mem[1297] = 4'b0000;
	mem[1298] = 4'b0000;
	mem[1299] = 4'b0000;
	mem[1300] = 4'b0000;
	mem[1301] = 4'b0000;
	mem[1302] = 4'b0000;
	mem[1303] = 4'b0000;
	mem[1304] = 4'b0000;
	mem[1305] = 4'b0000;
	mem[1306] = 4'b0000;
	mem[1307] = 4'b0000;
	mem[1308] = 4'b0000;
	mem[1309] = 4'b0000;
	mem[1310] = 4'b0000;
	mem[1311] = 4'b0000;
	mem[1312] = 4'b0000;
	mem[1313] = 4'b0000;
	mem[1314] = 4'b0000;
	mem[1315] = 4'b0000;
	mem[1316] = 4'b0000;
	mem[1317] = 4'b0000;
	mem[1318] = 4'b0000;
	mem[1319] = 4'b0000;
	mem[1320] = 4'b0000;
	mem[1321] = 4'b0000;
	mem[1322] = 4'b0000;
	mem[1323] = 4'b0000;
	mem[1324] = 4'b0000;
	mem[1325] = 4'b0000;
	mem[1326] = 4'b0000;
	mem[1327] = 4'b0000;
	mem[1328] = 4'b0000;
	mem[1329] = 4'b0000;
	mem[1330] = 4'b0000;
	mem[1331] = 4'b0000;
	mem[1332] = 4'b0000;
	mem[1333] = 4'b0000;
	mem[1334] = 4'b0000;
	mem[1335] = 4'b0000;
	mem[1336] = 4'b0000;
	mem[1337] = 4'b0000;
	mem[1338] = 4'b0000;
	mem[1339] = 4'b0000;
	mem[1340] = 4'b0000;
	mem[1341] = 4'b0000;
	mem[1342] = 4'b0000;
	mem[1343] = 4'b0000;
	mem[1344] = 4'b0001;
	mem[1345] = 4'b0000;
	mem[1346] = 4'b0000;
	mem[1347] = 4'b0000;
	mem[1348] = 4'b0000;
	mem[1349] = 4'b0000;
	mem[1350] = 4'b0000;
	mem[1351] = 4'b0000;
	mem[1352] = 4'b0000;
	mem[1353] = 4'b0000;
	mem[1354] = 4'b0000;
	mem[1355] = 4'b0000;
	mem[1356] = 4'b0000;
	mem[1357] = 4'b0000;
	mem[1358] = 4'b0000;
	mem[1359] = 4'b0000;
	mem[1360] = 4'b0000;
	mem[1361] = 4'b0000;
	mem[1362] = 4'b0000;
	mem[1363] = 4'b0000;
	mem[1364] = 4'b0000;
	mem[1365] = 4'b0000;
	mem[1366] = 4'b0000;
	mem[1367] = 4'b0000;
	mem[1368] = 4'b0000;
	mem[1369] = 4'b0000;
	mem[1370] = 4'b0000;
	mem[1371] = 4'b0000;
	mem[1372] = 4'b0000;
	mem[1373] = 4'b0000;
	mem[1374] = 4'b0000;
	mem[1375] = 4'b0000;
	mem[1376] = 4'b0000;
	mem[1377] = 4'b0000;
	mem[1378] = 4'b0000;
	mem[1379] = 4'b0000;
	mem[1380] = 4'b0000;
	mem[1381] = 4'b0000;
	mem[1382] = 4'b0000;
	mem[1383] = 4'b0000;
	mem[1384] = 4'b0000;
	mem[1385] = 4'b0000;
	mem[1386] = 4'b0000;
	mem[1387] = 4'b0000;
	mem[1388] = 4'b0000;
	mem[1389] = 4'b0000;
	mem[1390] = 4'b0000;
	mem[1391] = 4'b0000;
	mem[1392] = 4'b0000;
	mem[1393] = 4'b0000;
	mem[1394] = 4'b0000;
	mem[1395] = 4'b0000;
	mem[1396] = 4'b0000;
	mem[1397] = 4'b0000;
	mem[1398] = 4'b0000;
	mem[1399] = 4'b0000;
	mem[1400] = 4'b0000;
	mem[1401] = 4'b0000;
	mem[1402] = 4'b0000;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0101;
	mem[1412] = 4'b0111;
	mem[1413] = 4'b0111;
	mem[1414] = 4'b0111;
	mem[1415] = 4'b0111;
	mem[1416] = 4'b0111;
	mem[1417] = 4'b0111;
	mem[1418] = 4'b0111;
	mem[1419] = 4'b0111;
	mem[1420] = 4'b0111;
	mem[1421] = 4'b0111;
	mem[1422] = 4'b0111;
	mem[1423] = 4'b0111;
	mem[1424] = 4'b0111;
	mem[1425] = 4'b0111;
	mem[1426] = 4'b0111;
	mem[1427] = 4'b0111;
	mem[1428] = 4'b0010;
	mem[1429] = 4'b0000;
	mem[1430] = 4'b0000;
	mem[1431] = 4'b0000;
	mem[1432] = 4'b0000;
	mem[1433] = 4'b0000;
	mem[1434] = 4'b0000;
	mem[1435] = 4'b0000;
	mem[1436] = 4'b0000;
	mem[1437] = 4'b0000;
	mem[1438] = 4'b0000;
	mem[1439] = 4'b0000;
	mem[1440] = 4'b0000;
	mem[1441] = 4'b0000;
	mem[1442] = 4'b0000;
	mem[1443] = 4'b0000;
	mem[1444] = 4'b0000;
	mem[1445] = 4'b0111;
	mem[1446] = 4'b1001;
	mem[1447] = 4'b1001;
	mem[1448] = 4'b1001;
	mem[1449] = 4'b1001;
	mem[1450] = 4'b1001;
	mem[1451] = 4'b1001;
	mem[1452] = 4'b1001;
	mem[1453] = 4'b1001;
	mem[1454] = 4'b1001;
	mem[1455] = 4'b1001;
	mem[1456] = 4'b1001;
	mem[1457] = 4'b1001;
	mem[1458] = 4'b1001;
	mem[1459] = 4'b1001;
	mem[1460] = 4'b1001;
	mem[1461] = 4'b1001;
	mem[1462] = 4'b0011;
	mem[1463] = 4'b0000;
	mem[1464] = 4'b0000;
	mem[1465] = 4'b0000;
	mem[1466] = 4'b0000;
	mem[1467] = 4'b0000;
	mem[1468] = 4'b0000;
	mem[1469] = 4'b0000;
	mem[1470] = 4'b0000;
	mem[1471] = 4'b0000;
	mem[1472] = 4'b0000;
	mem[1473] = 4'b0000;
	mem[1474] = 4'b0000;
	mem[1475] = 4'b0000;
	mem[1476] = 4'b0000;
	mem[1477] = 4'b0000;
	mem[1478] = 4'b0000;
	mem[1479] = 4'b0110;
	mem[1480] = 4'b1001;
	mem[1481] = 4'b1010;
	mem[1482] = 4'b1001;
	mem[1483] = 4'b1001;
	mem[1484] = 4'b1001;
	mem[1485] = 4'b1001;
	mem[1486] = 4'b1001;
	mem[1487] = 4'b1001;
	mem[1488] = 4'b1001;
	mem[1489] = 4'b1001;
	mem[1490] = 4'b1001;
	mem[1491] = 4'b1001;
	mem[1492] = 4'b1001;
	mem[1493] = 4'b1001;
	mem[1494] = 4'b1001;
	mem[1495] = 4'b1001;
	mem[1496] = 4'b0010;
	mem[1497] = 4'b0000;
	mem[1498] = 4'b0000;
	mem[1499] = 4'b0000;
	mem[1500] = 4'b0000;
	mem[1501] = 4'b0000;
	mem[1502] = 4'b0000;
	mem[1503] = 4'b0000;
	mem[1504] = 4'b0000;
	mem[1505] = 4'b0000;
	mem[1506] = 4'b0000;
	mem[1507] = 4'b0000;
	mem[1508] = 4'b0000;
	mem[1509] = 4'b0000;
	mem[1510] = 4'b0000;
	mem[1511] = 4'b0000;
	mem[1512] = 4'b0000;
	mem[1513] = 4'b0110;
	mem[1514] = 4'b1001;
	mem[1515] = 4'b1001;
	mem[1516] = 4'b1000;
	mem[1517] = 4'b1000;
	mem[1518] = 4'b1000;
	mem[1519] = 4'b1000;
	mem[1520] = 4'b1000;
	mem[1521] = 4'b1000;
	mem[1522] = 4'b1000;
	mem[1523] = 4'b1000;
	mem[1524] = 4'b1000;
	mem[1525] = 4'b1001;
	mem[1526] = 4'b1001;
	mem[1527] = 4'b1001;
	mem[1528] = 4'b1001;
	mem[1529] = 4'b1001;
	mem[1530] = 4'b0001;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0111;
	mem[1540] = 4'b1100;
	mem[1541] = 4'b1100;
	mem[1542] = 4'b1100;
	mem[1543] = 4'b1100;
	mem[1544] = 4'b1100;
	mem[1545] = 4'b1100;
	mem[1546] = 4'b1100;
	mem[1547] = 4'b1100;
	mem[1548] = 4'b1100;
	mem[1549] = 4'b1100;
	mem[1550] = 4'b1100;
	mem[1551] = 4'b1100;
	mem[1552] = 4'b1100;
	mem[1553] = 4'b1100;
	mem[1554] = 4'b1100;
	mem[1555] = 4'b1100;
	mem[1556] = 4'b0011;
	mem[1557] = 4'b0000;
	mem[1558] = 4'b0000;
	mem[1559] = 4'b0000;
	mem[1560] = 4'b0000;
	mem[1561] = 4'b0000;
	mem[1562] = 4'b0000;
	mem[1563] = 4'b0000;
	mem[1564] = 4'b0000;
	mem[1565] = 4'b0000;
	mem[1566] = 4'b0000;
	mem[1567] = 4'b0000;
	mem[1568] = 4'b0000;
	mem[1569] = 4'b0000;
	mem[1570] = 4'b0000;
	mem[1571] = 4'b0000;
	mem[1572] = 4'b0000;
	mem[1573] = 4'b1100;
	mem[1574] = 4'b1111;
	mem[1575] = 4'b1111;
	mem[1576] = 4'b1111;
	mem[1577] = 4'b1111;
	mem[1578] = 4'b1111;
	mem[1579] = 4'b1111;
	mem[1580] = 4'b1111;
	mem[1581] = 4'b1111;
	mem[1582] = 4'b1111;
	mem[1583] = 4'b1111;
	mem[1584] = 4'b1111;
	mem[1585] = 4'b1111;
	mem[1586] = 4'b1111;
	mem[1587] = 4'b1111;
	mem[1588] = 4'b1111;
	mem[1589] = 4'b1111;
	mem[1590] = 4'b0110;
	mem[1591] = 4'b0000;
	mem[1592] = 4'b0000;
	mem[1593] = 4'b0000;
	mem[1594] = 4'b0000;
	mem[1595] = 4'b0000;
	mem[1596] = 4'b0000;
	mem[1597] = 4'b0000;
	mem[1598] = 4'b0000;
	mem[1599] = 4'b0000;
	mem[1600] = 4'b0000;
	mem[1601] = 4'b0000;
	mem[1602] = 4'b0000;
	mem[1603] = 4'b0000;
	mem[1604] = 4'b0000;
	mem[1605] = 4'b0000;
	mem[1606] = 4'b0001;
	mem[1607] = 4'b1100;
	mem[1608] = 4'b1111;
	mem[1609] = 4'b1111;
	mem[1610] = 4'b1111;
	mem[1611] = 4'b1111;
	mem[1612] = 4'b1111;
	mem[1613] = 4'b1111;
	mem[1614] = 4'b1111;
	mem[1615] = 4'b1111;
	mem[1616] = 4'b1111;
	mem[1617] = 4'b1111;
	mem[1618] = 4'b1111;
	mem[1619] = 4'b1111;
	mem[1620] = 4'b1111;
	mem[1621] = 4'b1111;
	mem[1622] = 4'b1111;
	mem[1623] = 4'b1111;
	mem[1624] = 4'b0100;
	mem[1625] = 4'b0000;
	mem[1626] = 4'b0000;
	mem[1627] = 4'b0000;
	mem[1628] = 4'b0000;
	mem[1629] = 4'b0000;
	mem[1630] = 4'b0000;
	mem[1631] = 4'b0000;
	mem[1632] = 4'b0000;
	mem[1633] = 4'b0000;
	mem[1634] = 4'b0000;
	mem[1635] = 4'b0000;
	mem[1636] = 4'b0000;
	mem[1637] = 4'b0000;
	mem[1638] = 4'b0000;
	mem[1639] = 4'b0000;
	mem[1640] = 4'b0000;
	mem[1641] = 4'b1001;
	mem[1642] = 4'b1110;
	mem[1643] = 4'b1101;
	mem[1644] = 4'b1101;
	mem[1645] = 4'b1101;
	mem[1646] = 4'b1110;
	mem[1647] = 4'b1110;
	mem[1648] = 4'b1110;
	mem[1649] = 4'b1101;
	mem[1650] = 4'b1101;
	mem[1651] = 4'b1101;
	mem[1652] = 4'b1101;
	mem[1653] = 4'b1101;
	mem[1654] = 4'b1111;
	mem[1655] = 4'b1111;
	mem[1656] = 4'b1111;
	mem[1657] = 4'b1111;
	mem[1658] = 4'b0010;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0111;
	mem[1668] = 4'b1100;
	mem[1669] = 4'b1101;
	mem[1670] = 4'b1101;
	mem[1671] = 4'b1101;
	mem[1672] = 4'b1101;
	mem[1673] = 4'b1101;
	mem[1674] = 4'b1101;
	mem[1675] = 4'b1101;
	mem[1676] = 4'b1101;
	mem[1677] = 4'b1101;
	mem[1678] = 4'b1101;
	mem[1679] = 4'b1101;
	mem[1680] = 4'b1101;
	mem[1681] = 4'b1101;
	mem[1682] = 4'b1101;
	mem[1683] = 4'b1101;
	mem[1684] = 4'b0110;
	mem[1685] = 4'b0100;
	mem[1686] = 4'b0100;
	mem[1687] = 4'b0100;
	mem[1688] = 4'b0100;
	mem[1689] = 4'b0100;
	mem[1690] = 4'b0100;
	mem[1691] = 4'b0100;
	mem[1692] = 4'b0100;
	mem[1693] = 4'b0100;
	mem[1694] = 4'b0100;
	mem[1695] = 4'b0100;
	mem[1696] = 4'b0100;
	mem[1697] = 4'b0100;
	mem[1698] = 4'b0100;
	mem[1699] = 4'b0100;
	mem[1700] = 4'b0100;
	mem[1701] = 4'b1101;
	mem[1702] = 4'b1111;
	mem[1703] = 4'b1111;
	mem[1704] = 4'b1111;
	mem[1705] = 4'b1111;
	mem[1706] = 4'b1111;
	mem[1707] = 4'b1111;
	mem[1708] = 4'b1111;
	mem[1709] = 4'b1111;
	mem[1710] = 4'b1111;
	mem[1711] = 4'b1111;
	mem[1712] = 4'b1111;
	mem[1713] = 4'b1111;
	mem[1714] = 4'b1111;
	mem[1715] = 4'b1111;
	mem[1716] = 4'b1111;
	mem[1717] = 4'b1111;
	mem[1718] = 4'b1001;
	mem[1719] = 4'b0100;
	mem[1720] = 4'b0100;
	mem[1721] = 4'b0100;
	mem[1722] = 4'b0100;
	mem[1723] = 4'b0100;
	mem[1724] = 4'b0101;
	mem[1725] = 4'b0101;
	mem[1726] = 4'b0101;
	mem[1727] = 4'b0101;
	mem[1728] = 4'b0100;
	mem[1729] = 4'b0100;
	mem[1730] = 4'b0100;
	mem[1731] = 4'b0101;
	mem[1732] = 4'b0100;
	mem[1733] = 4'b0100;
	mem[1734] = 4'b0101;
	mem[1735] = 4'b1101;
	mem[1736] = 4'b1111;
	mem[1737] = 4'b1111;
	mem[1738] = 4'b1111;
	mem[1739] = 4'b1111;
	mem[1740] = 4'b1111;
	mem[1741] = 4'b1111;
	mem[1742] = 4'b1111;
	mem[1743] = 4'b1111;
	mem[1744] = 4'b1111;
	mem[1745] = 4'b1111;
	mem[1746] = 4'b1111;
	mem[1747] = 4'b1111;
	mem[1748] = 4'b1111;
	mem[1749] = 4'b1111;
	mem[1750] = 4'b1111;
	mem[1751] = 4'b1111;
	mem[1752] = 4'b1000;
	mem[1753] = 4'b0101;
	mem[1754] = 4'b0101;
	mem[1755] = 4'b0101;
	mem[1756] = 4'b0101;
	mem[1757] = 4'b0101;
	mem[1758] = 4'b0101;
	mem[1759] = 4'b0101;
	mem[1760] = 4'b0101;
	mem[1761] = 4'b0101;
	mem[1762] = 4'b0101;
	mem[1763] = 4'b0101;
	mem[1764] = 4'b0101;
	mem[1765] = 4'b0101;
	mem[1766] = 4'b0101;
	mem[1767] = 4'b0101;
	mem[1768] = 4'b0101;
	mem[1769] = 4'b1011;
	mem[1770] = 4'b1101;
	mem[1771] = 4'b1101;
	mem[1772] = 4'b1101;
	mem[1773] = 4'b1110;
	mem[1774] = 4'b1111;
	mem[1775] = 4'b1111;
	mem[1776] = 4'b1111;
	mem[1777] = 4'b1111;
	mem[1778] = 4'b1101;
	mem[1779] = 4'b1101;
	mem[1780] = 4'b1101;
	mem[1781] = 4'b1101;
	mem[1782] = 4'b1101;
	mem[1783] = 4'b1111;
	mem[1784] = 4'b1111;
	mem[1785] = 4'b1111;
	mem[1786] = 4'b0010;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0111;
	mem[1796] = 4'b1100;
	mem[1797] = 4'b1101;
	mem[1798] = 4'b1101;
	mem[1799] = 4'b1101;
	mem[1800] = 4'b1101;
	mem[1801] = 4'b1101;
	mem[1802] = 4'b1101;
	mem[1803] = 4'b1101;
	mem[1804] = 4'b1101;
	mem[1805] = 4'b1101;
	mem[1806] = 4'b1101;
	mem[1807] = 4'b1101;
	mem[1808] = 4'b1101;
	mem[1809] = 4'b1101;
	mem[1810] = 4'b1101;
	mem[1811] = 4'b1101;
	mem[1812] = 4'b0110;
	mem[1813] = 4'b0100;
	mem[1814] = 4'b0100;
	mem[1815] = 4'b0100;
	mem[1816] = 4'b0100;
	mem[1817] = 4'b0100;
	mem[1818] = 4'b0100;
	mem[1819] = 4'b0100;
	mem[1820] = 4'b0100;
	mem[1821] = 4'b0100;
	mem[1822] = 4'b0100;
	mem[1823] = 4'b0100;
	mem[1824] = 4'b0100;
	mem[1825] = 4'b0101;
	mem[1826] = 4'b0101;
	mem[1827] = 4'b0101;
	mem[1828] = 4'b0101;
	mem[1829] = 4'b1101;
	mem[1830] = 4'b1111;
	mem[1831] = 4'b1111;
	mem[1832] = 4'b1111;
	mem[1833] = 4'b1111;
	mem[1834] = 4'b1111;
	mem[1835] = 4'b1111;
	mem[1836] = 4'b1111;
	mem[1837] = 4'b1111;
	mem[1838] = 4'b1111;
	mem[1839] = 4'b1111;
	mem[1840] = 4'b1111;
	mem[1841] = 4'b1111;
	mem[1842] = 4'b1111;
	mem[1843] = 4'b1111;
	mem[1844] = 4'b1111;
	mem[1845] = 4'b1111;
	mem[1846] = 4'b1001;
	mem[1847] = 4'b0101;
	mem[1848] = 4'b0101;
	mem[1849] = 4'b0101;
	mem[1850] = 4'b0101;
	mem[1851] = 4'b0101;
	mem[1852] = 4'b0101;
	mem[1853] = 4'b0101;
	mem[1854] = 4'b0101;
	mem[1855] = 4'b0101;
	mem[1856] = 4'b0110;
	mem[1857] = 4'b0101;
	mem[1858] = 4'b0101;
	mem[1859] = 4'b0101;
	mem[1860] = 4'b0101;
	mem[1861] = 4'b0110;
	mem[1862] = 4'b0110;
	mem[1863] = 4'b1101;
	mem[1864] = 4'b1111;
	mem[1865] = 4'b1111;
	mem[1866] = 4'b1111;
	mem[1867] = 4'b1111;
	mem[1868] = 4'b1111;
	mem[1869] = 4'b1111;
	mem[1870] = 4'b1111;
	mem[1871] = 4'b1111;
	mem[1872] = 4'b1111;
	mem[1873] = 4'b1111;
	mem[1874] = 4'b1111;
	mem[1875] = 4'b1111;
	mem[1876] = 4'b1111;
	mem[1877] = 4'b1111;
	mem[1878] = 4'b1111;
	mem[1879] = 4'b1111;
	mem[1880] = 4'b1000;
	mem[1881] = 4'b0110;
	mem[1882] = 4'b0110;
	mem[1883] = 4'b0110;
	mem[1884] = 4'b0110;
	mem[1885] = 4'b0110;
	mem[1886] = 4'b0110;
	mem[1887] = 4'b0110;
	mem[1888] = 4'b0110;
	mem[1889] = 4'b0110;
	mem[1890] = 4'b0110;
	mem[1891] = 4'b0110;
	mem[1892] = 4'b0110;
	mem[1893] = 4'b0110;
	mem[1894] = 4'b0110;
	mem[1895] = 4'b0110;
	mem[1896] = 4'b0110;
	mem[1897] = 4'b1011;
	mem[1898] = 4'b1101;
	mem[1899] = 4'b1101;
	mem[1900] = 4'b1110;
	mem[1901] = 4'b1111;
	mem[1902] = 4'b1111;
	mem[1903] = 4'b1111;
	mem[1904] = 4'b1111;
	mem[1905] = 4'b1111;
	mem[1906] = 4'b1111;
	mem[1907] = 4'b1101;
	mem[1908] = 4'b1101;
	mem[1909] = 4'b1101;
	mem[1910] = 4'b1101;
	mem[1911] = 4'b1101;
	mem[1912] = 4'b1111;
	mem[1913] = 4'b1111;
	mem[1914] = 4'b0011;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0111;
	mem[1924] = 4'b1100;
	mem[1925] = 4'b1101;
	mem[1926] = 4'b1101;
	mem[1927] = 4'b1101;
	mem[1928] = 4'b1101;
	mem[1929] = 4'b1101;
	mem[1930] = 4'b1101;
	mem[1931] = 4'b1101;
	mem[1932] = 4'b1101;
	mem[1933] = 4'b1101;
	mem[1934] = 4'b1101;
	mem[1935] = 4'b1101;
	mem[1936] = 4'b1101;
	mem[1937] = 4'b1101;
	mem[1938] = 4'b1101;
	mem[1939] = 4'b1101;
	mem[1940] = 4'b0110;
	mem[1941] = 4'b0100;
	mem[1942] = 4'b0100;
	mem[1943] = 4'b0100;
	mem[1944] = 4'b0100;
	mem[1945] = 4'b0100;
	mem[1946] = 4'b0100;
	mem[1947] = 4'b0100;
	mem[1948] = 4'b0100;
	mem[1949] = 4'b0100;
	mem[1950] = 4'b0100;
	mem[1951] = 4'b0101;
	mem[1952] = 4'b0101;
	mem[1953] = 4'b0101;
	mem[1954] = 4'b0101;
	mem[1955] = 4'b0101;
	mem[1956] = 4'b0101;
	mem[1957] = 4'b1101;
	mem[1958] = 4'b1111;
	mem[1959] = 4'b1111;
	mem[1960] = 4'b1111;
	mem[1961] = 4'b1111;
	mem[1962] = 4'b1111;
	mem[1963] = 4'b1111;
	mem[1964] = 4'b1111;
	mem[1965] = 4'b1111;
	mem[1966] = 4'b1111;
	mem[1967] = 4'b1111;
	mem[1968] = 4'b1111;
	mem[1969] = 4'b1111;
	mem[1970] = 4'b1111;
	mem[1971] = 4'b1111;
	mem[1972] = 4'b1111;
	mem[1973] = 4'b1111;
	mem[1974] = 4'b1001;
	mem[1975] = 4'b0101;
	mem[1976] = 4'b0101;
	mem[1977] = 4'b0101;
	mem[1978] = 4'b0101;
	mem[1979] = 4'b0101;
	mem[1980] = 4'b0101;
	mem[1981] = 4'b0101;
	mem[1982] = 4'b0101;
	mem[1983] = 4'b0101;
	mem[1984] = 4'b0101;
	mem[1985] = 4'b0110;
	mem[1986] = 4'b0110;
	mem[1987] = 4'b0110;
	mem[1988] = 4'b0110;
	mem[1989] = 4'b0110;
	mem[1990] = 4'b0110;
	mem[1991] = 4'b1101;
	mem[1992] = 4'b1111;
	mem[1993] = 4'b1111;
	mem[1994] = 4'b1111;
	mem[1995] = 4'b1111;
	mem[1996] = 4'b1111;
	mem[1997] = 4'b1111;
	mem[1998] = 4'b1111;
	mem[1999] = 4'b1111;
	mem[2000] = 4'b1111;
	mem[2001] = 4'b1111;
	mem[2002] = 4'b1111;
	mem[2003] = 4'b1111;
	mem[2004] = 4'b1111;
	mem[2005] = 4'b1111;
	mem[2006] = 4'b1111;
	mem[2007] = 4'b1111;
	mem[2008] = 4'b1000;
	mem[2009] = 4'b0110;
	mem[2010] = 4'b0110;
	mem[2011] = 4'b0110;
	mem[2012] = 4'b0110;
	mem[2013] = 4'b0110;
	mem[2014] = 4'b0110;
	mem[2015] = 4'b0110;
	mem[2016] = 4'b0110;
	mem[2017] = 4'b0110;
	mem[2018] = 4'b0110;
	mem[2019] = 4'b0110;
	mem[2020] = 4'b0110;
	mem[2021] = 4'b0110;
	mem[2022] = 4'b0110;
	mem[2023] = 4'b0110;
	mem[2024] = 4'b0110;
	mem[2025] = 4'b1011;
	mem[2026] = 4'b1101;
	mem[2027] = 4'b1101;
	mem[2028] = 4'b1111;
	mem[2029] = 4'b1111;
	mem[2030] = 4'b1111;
	mem[2031] = 4'b1111;
	mem[2032] = 4'b1111;
	mem[2033] = 4'b1111;
	mem[2034] = 4'b1111;
	mem[2035] = 4'b1111;
	mem[2036] = 4'b1101;
	mem[2037] = 4'b1101;
	mem[2038] = 4'b1101;
	mem[2039] = 4'b1101;
	mem[2040] = 4'b1101;
	mem[2041] = 4'b1110;
	mem[2042] = 4'b0011;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0111;
	mem[2052] = 4'b1100;
	mem[2053] = 4'b1101;
	mem[2054] = 4'b1101;
	mem[2055] = 4'b1101;
	mem[2056] = 4'b1101;
	mem[2057] = 4'b1101;
	mem[2058] = 4'b1101;
	mem[2059] = 4'b1101;
	mem[2060] = 4'b1101;
	mem[2061] = 4'b1101;
	mem[2062] = 4'b1101;
	mem[2063] = 4'b1101;
	mem[2064] = 4'b1101;
	mem[2065] = 4'b1101;
	mem[2066] = 4'b1101;
	mem[2067] = 4'b1101;
	mem[2068] = 4'b0111;
	mem[2069] = 4'b0100;
	mem[2070] = 4'b0100;
	mem[2071] = 4'b0100;
	mem[2072] = 4'b0100;
	mem[2073] = 4'b0100;
	mem[2074] = 4'b0100;
	mem[2075] = 4'b0100;
	mem[2076] = 4'b0100;
	mem[2077] = 4'b0101;
	mem[2078] = 4'b0101;
	mem[2079] = 4'b0101;
	mem[2080] = 4'b0101;
	mem[2081] = 4'b0101;
	mem[2082] = 4'b0101;
	mem[2083] = 4'b0101;
	mem[2084] = 4'b0101;
	mem[2085] = 4'b1101;
	mem[2086] = 4'b1111;
	mem[2087] = 4'b1111;
	mem[2088] = 4'b1111;
	mem[2089] = 4'b1111;
	mem[2090] = 4'b1111;
	mem[2091] = 4'b1111;
	mem[2092] = 4'b1111;
	mem[2093] = 4'b1111;
	mem[2094] = 4'b1111;
	mem[2095] = 4'b1111;
	mem[2096] = 4'b1111;
	mem[2097] = 4'b1111;
	mem[2098] = 4'b1111;
	mem[2099] = 4'b1111;
	mem[2100] = 4'b1111;
	mem[2101] = 4'b1111;
	mem[2102] = 4'b1001;
	mem[2103] = 4'b0101;
	mem[2104] = 4'b0101;
	mem[2105] = 4'b0101;
	mem[2106] = 4'b0110;
	mem[2107] = 4'b0110;
	mem[2108] = 4'b0110;
	mem[2109] = 4'b0101;
	mem[2110] = 4'b0101;
	mem[2111] = 4'b0101;
	mem[2112] = 4'b0110;
	mem[2113] = 4'b0101;
	mem[2114] = 4'b0110;
	mem[2115] = 4'b0110;
	mem[2116] = 4'b0110;
	mem[2117] = 4'b0110;
	mem[2118] = 4'b0110;
	mem[2119] = 4'b1101;
	mem[2120] = 4'b1111;
	mem[2121] = 4'b1111;
	mem[2122] = 4'b1111;
	mem[2123] = 4'b1111;
	mem[2124] = 4'b1111;
	mem[2125] = 4'b1111;
	mem[2126] = 4'b1111;
	mem[2127] = 4'b1111;
	mem[2128] = 4'b1111;
	mem[2129] = 4'b1111;
	mem[2130] = 4'b1111;
	mem[2131] = 4'b1111;
	mem[2132] = 4'b1111;
	mem[2133] = 4'b1111;
	mem[2134] = 4'b1111;
	mem[2135] = 4'b1111;
	mem[2136] = 4'b1000;
	mem[2137] = 4'b0110;
	mem[2138] = 4'b0110;
	mem[2139] = 4'b0110;
	mem[2140] = 4'b0110;
	mem[2141] = 4'b0110;
	mem[2142] = 4'b0110;
	mem[2143] = 4'b0110;
	mem[2144] = 4'b0110;
	mem[2145] = 4'b0110;
	mem[2146] = 4'b0110;
	mem[2147] = 4'b0110;
	mem[2148] = 4'b0110;
	mem[2149] = 4'b0110;
	mem[2150] = 4'b0110;
	mem[2151] = 4'b0110;
	mem[2152] = 4'b0110;
	mem[2153] = 4'b1011;
	mem[2154] = 4'b1101;
	mem[2155] = 4'b1101;
	mem[2156] = 4'b1111;
	mem[2157] = 4'b1111;
	mem[2158] = 4'b1111;
	mem[2159] = 4'b1111;
	mem[2160] = 4'b1111;
	mem[2161] = 4'b1111;
	mem[2162] = 4'b1111;
	mem[2163] = 4'b1111;
	mem[2164] = 4'b1111;
	mem[2165] = 4'b1101;
	mem[2166] = 4'b1101;
	mem[2167] = 4'b1101;
	mem[2168] = 4'b1101;
	mem[2169] = 4'b1101;
	mem[2170] = 4'b0100;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0111;
	mem[2180] = 4'b1100;
	mem[2181] = 4'b1101;
	mem[2182] = 4'b1101;
	mem[2183] = 4'b1101;
	mem[2184] = 4'b1101;
	mem[2185] = 4'b1101;
	mem[2186] = 4'b1101;
	mem[2187] = 4'b1101;
	mem[2188] = 4'b1101;
	mem[2189] = 4'b1101;
	mem[2190] = 4'b1101;
	mem[2191] = 4'b1101;
	mem[2192] = 4'b1101;
	mem[2193] = 4'b1101;
	mem[2194] = 4'b1101;
	mem[2195] = 4'b1101;
	mem[2196] = 4'b0111;
	mem[2197] = 4'b0100;
	mem[2198] = 4'b0100;
	mem[2199] = 4'b0100;
	mem[2200] = 4'b0100;
	mem[2201] = 4'b0100;
	mem[2202] = 4'b0100;
	mem[2203] = 4'b0100;
	mem[2204] = 4'b0101;
	mem[2205] = 4'b0101;
	mem[2206] = 4'b0101;
	mem[2207] = 4'b0101;
	mem[2208] = 4'b0101;
	mem[2209] = 4'b0101;
	mem[2210] = 4'b0101;
	mem[2211] = 4'b0101;
	mem[2212] = 4'b0101;
	mem[2213] = 4'b1101;
	mem[2214] = 4'b1111;
	mem[2215] = 4'b1111;
	mem[2216] = 4'b1111;
	mem[2217] = 4'b1111;
	mem[2218] = 4'b1111;
	mem[2219] = 4'b1111;
	mem[2220] = 4'b1111;
	mem[2221] = 4'b1111;
	mem[2222] = 4'b1111;
	mem[2223] = 4'b1111;
	mem[2224] = 4'b1111;
	mem[2225] = 4'b1111;
	mem[2226] = 4'b1111;
	mem[2227] = 4'b1111;
	mem[2228] = 4'b1111;
	mem[2229] = 4'b1111;
	mem[2230] = 4'b1000;
	mem[2231] = 4'b0101;
	mem[2232] = 4'b0101;
	mem[2233] = 4'b0110;
	mem[2234] = 4'b0110;
	mem[2235] = 4'b0101;
	mem[2236] = 4'b0101;
	mem[2237] = 4'b0110;
	mem[2238] = 4'b0101;
	mem[2239] = 4'b0101;
	mem[2240] = 4'b0110;
	mem[2241] = 4'b0110;
	mem[2242] = 4'b0101;
	mem[2243] = 4'b0101;
	mem[2244] = 4'b0110;
	mem[2245] = 4'b0110;
	mem[2246] = 4'b0110;
	mem[2247] = 4'b1101;
	mem[2248] = 4'b1111;
	mem[2249] = 4'b1111;
	mem[2250] = 4'b1111;
	mem[2251] = 4'b1111;
	mem[2252] = 4'b1111;
	mem[2253] = 4'b1111;
	mem[2254] = 4'b1111;
	mem[2255] = 4'b1111;
	mem[2256] = 4'b1111;
	mem[2257] = 4'b1111;
	mem[2258] = 4'b1111;
	mem[2259] = 4'b1111;
	mem[2260] = 4'b1111;
	mem[2261] = 4'b1111;
	mem[2262] = 4'b1111;
	mem[2263] = 4'b1111;
	mem[2264] = 4'b1000;
	mem[2265] = 4'b0110;
	mem[2266] = 4'b0110;
	mem[2267] = 4'b0110;
	mem[2268] = 4'b0110;
	mem[2269] = 4'b0110;
	mem[2270] = 4'b0110;
	mem[2271] = 4'b0110;
	mem[2272] = 4'b0110;
	mem[2273] = 4'b0110;
	mem[2274] = 4'b0110;
	mem[2275] = 4'b0110;
	mem[2276] = 4'b0110;
	mem[2277] = 4'b0110;
	mem[2278] = 4'b0110;
	mem[2279] = 4'b0110;
	mem[2280] = 4'b0110;
	mem[2281] = 4'b1011;
	mem[2282] = 4'b1101;
	mem[2283] = 4'b1101;
	mem[2284] = 4'b1110;
	mem[2285] = 4'b1111;
	mem[2286] = 4'b1111;
	mem[2287] = 4'b1111;
	mem[2288] = 4'b1111;
	mem[2289] = 4'b1111;
	mem[2290] = 4'b1111;
	mem[2291] = 4'b1111;
	mem[2292] = 4'b1111;
	mem[2293] = 4'b1101;
	mem[2294] = 4'b1101;
	mem[2295] = 4'b1101;
	mem[2296] = 4'b1101;
	mem[2297] = 4'b1101;
	mem[2298] = 4'b0011;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0111;
	mem[2308] = 4'b1100;
	mem[2309] = 4'b1101;
	mem[2310] = 4'b1101;
	mem[2311] = 4'b1101;
	mem[2312] = 4'b1101;
	mem[2313] = 4'b1101;
	mem[2314] = 4'b1101;
	mem[2315] = 4'b1101;
	mem[2316] = 4'b1101;
	mem[2317] = 4'b1101;
	mem[2318] = 4'b1101;
	mem[2319] = 4'b1101;
	mem[2320] = 4'b1101;
	mem[2321] = 4'b1101;
	mem[2322] = 4'b1101;
	mem[2323] = 4'b1101;
	mem[2324] = 4'b0111;
	mem[2325] = 4'b0100;
	mem[2326] = 4'b0100;
	mem[2327] = 4'b0100;
	mem[2328] = 4'b0100;
	mem[2329] = 4'b0100;
	mem[2330] = 4'b0101;
	mem[2331] = 4'b0101;
	mem[2332] = 4'b0101;
	mem[2333] = 4'b0101;
	mem[2334] = 4'b0101;
	mem[2335] = 4'b0101;
	mem[2336] = 4'b0101;
	mem[2337] = 4'b0101;
	mem[2338] = 4'b0101;
	mem[2339] = 4'b0101;
	mem[2340] = 4'b0101;
	mem[2341] = 4'b1101;
	mem[2342] = 4'b1111;
	mem[2343] = 4'b1111;
	mem[2344] = 4'b1111;
	mem[2345] = 4'b1111;
	mem[2346] = 4'b1111;
	mem[2347] = 4'b1111;
	mem[2348] = 4'b1111;
	mem[2349] = 4'b1111;
	mem[2350] = 4'b1111;
	mem[2351] = 4'b1111;
	mem[2352] = 4'b1111;
	mem[2353] = 4'b1111;
	mem[2354] = 4'b1111;
	mem[2355] = 4'b1111;
	mem[2356] = 4'b1111;
	mem[2357] = 4'b1111;
	mem[2358] = 4'b1001;
	mem[2359] = 4'b0101;
	mem[2360] = 4'b0101;
	mem[2361] = 4'b0101;
	mem[2362] = 4'b0110;
	mem[2363] = 4'b0101;
	mem[2364] = 4'b0101;
	mem[2365] = 4'b0101;
	mem[2366] = 4'b0110;
	mem[2367] = 4'b0101;
	mem[2368] = 4'b0101;
	mem[2369] = 4'b0110;
	mem[2370] = 4'b0110;
	mem[2371] = 4'b0110;
	mem[2372] = 4'b0110;
	mem[2373] = 4'b0110;
	mem[2374] = 4'b0110;
	mem[2375] = 4'b1101;
	mem[2376] = 4'b1111;
	mem[2377] = 4'b1111;
	mem[2378] = 4'b1111;
	mem[2379] = 4'b1111;
	mem[2380] = 4'b1111;
	mem[2381] = 4'b1111;
	mem[2382] = 4'b1111;
	mem[2383] = 4'b1111;
	mem[2384] = 4'b1111;
	mem[2385] = 4'b1111;
	mem[2386] = 4'b1111;
	mem[2387] = 4'b1111;
	mem[2388] = 4'b1111;
	mem[2389] = 4'b1111;
	mem[2390] = 4'b1111;
	mem[2391] = 4'b1111;
	mem[2392] = 4'b1000;
	mem[2393] = 4'b0110;
	mem[2394] = 4'b0110;
	mem[2395] = 4'b0110;
	mem[2396] = 4'b0110;
	mem[2397] = 4'b0110;
	mem[2398] = 4'b0110;
	mem[2399] = 4'b0110;
	mem[2400] = 4'b0110;
	mem[2401] = 4'b0110;
	mem[2402] = 4'b0110;
	mem[2403] = 4'b0110;
	mem[2404] = 4'b0110;
	mem[2405] = 4'b0110;
	mem[2406] = 4'b0110;
	mem[2407] = 4'b0110;
	mem[2408] = 4'b0110;
	mem[2409] = 4'b1011;
	mem[2410] = 4'b1101;
	mem[2411] = 4'b1101;
	mem[2412] = 4'b1101;
	mem[2413] = 4'b1111;
	mem[2414] = 4'b1111;
	mem[2415] = 4'b1111;
	mem[2416] = 4'b1111;
	mem[2417] = 4'b1111;
	mem[2418] = 4'b1111;
	mem[2419] = 4'b1111;
	mem[2420] = 4'b1111;
	mem[2421] = 4'b1110;
	mem[2422] = 4'b1101;
	mem[2423] = 4'b1110;
	mem[2424] = 4'b1101;
	mem[2425] = 4'b1101;
	mem[2426] = 4'b0100;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0111;
	mem[2436] = 4'b1100;
	mem[2437] = 4'b1101;
	mem[2438] = 4'b1101;
	mem[2439] = 4'b1101;
	mem[2440] = 4'b1101;
	mem[2441] = 4'b1101;
	mem[2442] = 4'b1101;
	mem[2443] = 4'b1101;
	mem[2444] = 4'b1101;
	mem[2445] = 4'b1101;
	mem[2446] = 4'b1101;
	mem[2447] = 4'b1101;
	mem[2448] = 4'b1101;
	mem[2449] = 4'b1101;
	mem[2450] = 4'b1101;
	mem[2451] = 4'b1101;
	mem[2452] = 4'b0111;
	mem[2453] = 4'b0100;
	mem[2454] = 4'b0100;
	mem[2455] = 4'b0100;
	mem[2456] = 4'b0101;
	mem[2457] = 4'b0101;
	mem[2458] = 4'b0101;
	mem[2459] = 4'b0101;
	mem[2460] = 4'b0101;
	mem[2461] = 4'b0101;
	mem[2462] = 4'b0101;
	mem[2463] = 4'b0101;
	mem[2464] = 4'b0101;
	mem[2465] = 4'b0101;
	mem[2466] = 4'b0101;
	mem[2467] = 4'b0101;
	mem[2468] = 4'b0101;
	mem[2469] = 4'b1101;
	mem[2470] = 4'b1111;
	mem[2471] = 4'b1111;
	mem[2472] = 4'b1111;
	mem[2473] = 4'b1111;
	mem[2474] = 4'b1111;
	mem[2475] = 4'b1111;
	mem[2476] = 4'b1111;
	mem[2477] = 4'b1111;
	mem[2478] = 4'b1111;
	mem[2479] = 4'b1111;
	mem[2480] = 4'b1111;
	mem[2481] = 4'b1111;
	mem[2482] = 4'b1111;
	mem[2483] = 4'b1111;
	mem[2484] = 4'b1111;
	mem[2485] = 4'b1111;
	mem[2486] = 4'b1001;
	mem[2487] = 4'b0110;
	mem[2488] = 4'b0101;
	mem[2489] = 4'b0101;
	mem[2490] = 4'b0101;
	mem[2491] = 4'b0110;
	mem[2492] = 4'b0101;
	mem[2493] = 4'b0101;
	mem[2494] = 4'b0110;
	mem[2495] = 4'b0110;
	mem[2496] = 4'b0110;
	mem[2497] = 4'b0110;
	mem[2498] = 4'b0110;
	mem[2499] = 4'b0110;
	mem[2500] = 4'b0110;
	mem[2501] = 4'b0110;
	mem[2502] = 4'b0110;
	mem[2503] = 4'b1101;
	mem[2504] = 4'b1111;
	mem[2505] = 4'b1111;
	mem[2506] = 4'b1111;
	mem[2507] = 4'b1111;
	mem[2508] = 4'b1111;
	mem[2509] = 4'b1111;
	mem[2510] = 4'b1111;
	mem[2511] = 4'b1111;
	mem[2512] = 4'b1111;
	mem[2513] = 4'b1111;
	mem[2514] = 4'b1111;
	mem[2515] = 4'b1111;
	mem[2516] = 4'b1111;
	mem[2517] = 4'b1111;
	mem[2518] = 4'b1111;
	mem[2519] = 4'b1111;
	mem[2520] = 4'b1000;
	mem[2521] = 4'b0110;
	mem[2522] = 4'b0110;
	mem[2523] = 4'b0110;
	mem[2524] = 4'b0110;
	mem[2525] = 4'b0110;
	mem[2526] = 4'b0110;
	mem[2527] = 4'b0110;
	mem[2528] = 4'b0110;
	mem[2529] = 4'b0110;
	mem[2530] = 4'b0110;
	mem[2531] = 4'b0110;
	mem[2532] = 4'b0110;
	mem[2533] = 4'b0110;
	mem[2534] = 4'b0110;
	mem[2535] = 4'b0110;
	mem[2536] = 4'b0110;
	mem[2537] = 4'b1011;
	mem[2538] = 4'b1101;
	mem[2539] = 4'b1101;
	mem[2540] = 4'b1101;
	mem[2541] = 4'b1101;
	mem[2542] = 4'b1111;
	mem[2543] = 4'b1111;
	mem[2544] = 4'b1111;
	mem[2545] = 4'b1111;
	mem[2546] = 4'b1111;
	mem[2547] = 4'b1111;
	mem[2548] = 4'b1111;
	mem[2549] = 4'b1101;
	mem[2550] = 4'b1101;
	mem[2551] = 4'b1111;
	mem[2552] = 4'b1110;
	mem[2553] = 4'b1111;
	mem[2554] = 4'b0100;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b0111;
	mem[2564] = 4'b1100;
	mem[2565] = 4'b1101;
	mem[2566] = 4'b1101;
	mem[2567] = 4'b1101;
	mem[2568] = 4'b1101;
	mem[2569] = 4'b1101;
	mem[2570] = 4'b1101;
	mem[2571] = 4'b1101;
	mem[2572] = 4'b1101;
	mem[2573] = 4'b1101;
	mem[2574] = 4'b1101;
	mem[2575] = 4'b1101;
	mem[2576] = 4'b1101;
	mem[2577] = 4'b1101;
	mem[2578] = 4'b1101;
	mem[2579] = 4'b1101;
	mem[2580] = 4'b0111;
	mem[2581] = 4'b0100;
	mem[2582] = 4'b0101;
	mem[2583] = 4'b0101;
	mem[2584] = 4'b0101;
	mem[2585] = 4'b0101;
	mem[2586] = 4'b0101;
	mem[2587] = 4'b0101;
	mem[2588] = 4'b0101;
	mem[2589] = 4'b0101;
	mem[2590] = 4'b0101;
	mem[2591] = 4'b0101;
	mem[2592] = 4'b0101;
	mem[2593] = 4'b0101;
	mem[2594] = 4'b0101;
	mem[2595] = 4'b0101;
	mem[2596] = 4'b0101;
	mem[2597] = 4'b1101;
	mem[2598] = 4'b1111;
	mem[2599] = 4'b1111;
	mem[2600] = 4'b1111;
	mem[2601] = 4'b1111;
	mem[2602] = 4'b1111;
	mem[2603] = 4'b1111;
	mem[2604] = 4'b1111;
	mem[2605] = 4'b1111;
	mem[2606] = 4'b1111;
	mem[2607] = 4'b1111;
	mem[2608] = 4'b1111;
	mem[2609] = 4'b1111;
	mem[2610] = 4'b1111;
	mem[2611] = 4'b1111;
	mem[2612] = 4'b1110;
	mem[2613] = 4'b1111;
	mem[2614] = 4'b1001;
	mem[2615] = 4'b0101;
	mem[2616] = 4'b0110;
	mem[2617] = 4'b0101;
	mem[2618] = 4'b0101;
	mem[2619] = 4'b0110;
	mem[2620] = 4'b0110;
	mem[2621] = 4'b0101;
	mem[2622] = 4'b0110;
	mem[2623] = 4'b0110;
	mem[2624] = 4'b0110;
	mem[2625] = 4'b0110;
	mem[2626] = 4'b0110;
	mem[2627] = 4'b0110;
	mem[2628] = 4'b0110;
	mem[2629] = 4'b0110;
	mem[2630] = 4'b0110;
	mem[2631] = 4'b1101;
	mem[2632] = 4'b1111;
	mem[2633] = 4'b1111;
	mem[2634] = 4'b1111;
	mem[2635] = 4'b1111;
	mem[2636] = 4'b1111;
	mem[2637] = 4'b1111;
	mem[2638] = 4'b1111;
	mem[2639] = 4'b1111;
	mem[2640] = 4'b1111;
	mem[2641] = 4'b1111;
	mem[2642] = 4'b1111;
	mem[2643] = 4'b1111;
	mem[2644] = 4'b1111;
	mem[2645] = 4'b1111;
	mem[2646] = 4'b1111;
	mem[2647] = 4'b1111;
	mem[2648] = 4'b1000;
	mem[2649] = 4'b0110;
	mem[2650] = 4'b0110;
	mem[2651] = 4'b0110;
	mem[2652] = 4'b0110;
	mem[2653] = 4'b0110;
	mem[2654] = 4'b0110;
	mem[2655] = 4'b0110;
	mem[2656] = 4'b0110;
	mem[2657] = 4'b0110;
	mem[2658] = 4'b0110;
	mem[2659] = 4'b0110;
	mem[2660] = 4'b0110;
	mem[2661] = 4'b0110;
	mem[2662] = 4'b0110;
	mem[2663] = 4'b0110;
	mem[2664] = 4'b0110;
	mem[2665] = 4'b1100;
	mem[2666] = 4'b1110;
	mem[2667] = 4'b1101;
	mem[2668] = 4'b1101;
	mem[2669] = 4'b1101;
	mem[2670] = 4'b1101;
	mem[2671] = 4'b1111;
	mem[2672] = 4'b1111;
	mem[2673] = 4'b1111;
	mem[2674] = 4'b1111;
	mem[2675] = 4'b1111;
	mem[2676] = 4'b1110;
	mem[2677] = 4'b1101;
	mem[2678] = 4'b1101;
	mem[2679] = 4'b1111;
	mem[2680] = 4'b1111;
	mem[2681] = 4'b1111;
	mem[2682] = 4'b0011;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b0111;
	mem[2692] = 4'b1100;
	mem[2693] = 4'b1101;
	mem[2694] = 4'b1101;
	mem[2695] = 4'b1101;
	mem[2696] = 4'b1101;
	mem[2697] = 4'b1101;
	mem[2698] = 4'b1101;
	mem[2699] = 4'b1101;
	mem[2700] = 4'b1101;
	mem[2701] = 4'b1101;
	mem[2702] = 4'b1101;
	mem[2703] = 4'b1101;
	mem[2704] = 4'b1101;
	mem[2705] = 4'b1101;
	mem[2706] = 4'b1101;
	mem[2707] = 4'b1101;
	mem[2708] = 4'b0111;
	mem[2709] = 4'b0101;
	mem[2710] = 4'b0101;
	mem[2711] = 4'b0101;
	mem[2712] = 4'b0101;
	mem[2713] = 4'b0101;
	mem[2714] = 4'b0101;
	mem[2715] = 4'b0101;
	mem[2716] = 4'b0101;
	mem[2717] = 4'b0101;
	mem[2718] = 4'b0101;
	mem[2719] = 4'b0101;
	mem[2720] = 4'b0101;
	mem[2721] = 4'b0101;
	mem[2722] = 4'b0101;
	mem[2723] = 4'b0101;
	mem[2724] = 4'b0101;
	mem[2725] = 4'b1101;
	mem[2726] = 4'b1111;
	mem[2727] = 4'b1111;
	mem[2728] = 4'b1111;
	mem[2729] = 4'b1111;
	mem[2730] = 4'b1111;
	mem[2731] = 4'b1111;
	mem[2732] = 4'b1111;
	mem[2733] = 4'b1111;
	mem[2734] = 4'b1111;
	mem[2735] = 4'b1111;
	mem[2736] = 4'b1111;
	mem[2737] = 4'b1111;
	mem[2738] = 4'b1110;
	mem[2739] = 4'b1101;
	mem[2740] = 4'b1101;
	mem[2741] = 4'b1101;
	mem[2742] = 4'b1001;
	mem[2743] = 4'b0101;
	mem[2744] = 4'b0101;
	mem[2745] = 4'b0110;
	mem[2746] = 4'b0101;
	mem[2747] = 4'b0101;
	mem[2748] = 4'b0110;
	mem[2749] = 4'b0110;
	mem[2750] = 4'b0110;
	mem[2751] = 4'b0110;
	mem[2752] = 4'b0110;
	mem[2753] = 4'b0110;
	mem[2754] = 4'b0110;
	mem[2755] = 4'b0110;
	mem[2756] = 4'b0110;
	mem[2757] = 4'b0110;
	mem[2758] = 4'b0110;
	mem[2759] = 4'b1101;
	mem[2760] = 4'b1111;
	mem[2761] = 4'b1111;
	mem[2762] = 4'b1111;
	mem[2763] = 4'b1111;
	mem[2764] = 4'b1111;
	mem[2765] = 4'b1111;
	mem[2766] = 4'b1111;
	mem[2767] = 4'b1111;
	mem[2768] = 4'b1111;
	mem[2769] = 4'b1111;
	mem[2770] = 4'b1111;
	mem[2771] = 4'b1111;
	mem[2772] = 4'b1111;
	mem[2773] = 4'b1111;
	mem[2774] = 4'b1111;
	mem[2775] = 4'b1111;
	mem[2776] = 4'b1001;
	mem[2777] = 4'b0110;
	mem[2778] = 4'b0110;
	mem[2779] = 4'b0110;
	mem[2780] = 4'b0110;
	mem[2781] = 4'b0110;
	mem[2782] = 4'b0110;
	mem[2783] = 4'b0110;
	mem[2784] = 4'b0110;
	mem[2785] = 4'b0110;
	mem[2786] = 4'b0110;
	mem[2787] = 4'b0110;
	mem[2788] = 4'b0110;
	mem[2789] = 4'b0111;
	mem[2790] = 4'b0111;
	mem[2791] = 4'b0110;
	mem[2792] = 4'b0111;
	mem[2793] = 4'b1100;
	mem[2794] = 4'b1111;
	mem[2795] = 4'b1101;
	mem[2796] = 4'b1101;
	mem[2797] = 4'b1101;
	mem[2798] = 4'b1101;
	mem[2799] = 4'b1101;
	mem[2800] = 4'b1110;
	mem[2801] = 4'b1110;
	mem[2802] = 4'b1110;
	mem[2803] = 4'b1110;
	mem[2804] = 4'b1101;
	mem[2805] = 4'b1101;
	mem[2806] = 4'b1110;
	mem[2807] = 4'b1111;
	mem[2808] = 4'b1111;
	mem[2809] = 4'b1111;
	mem[2810] = 4'b0011;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b0111;
	mem[2820] = 4'b1100;
	mem[2821] = 4'b1101;
	mem[2822] = 4'b1101;
	mem[2823] = 4'b1101;
	mem[2824] = 4'b1101;
	mem[2825] = 4'b1101;
	mem[2826] = 4'b1101;
	mem[2827] = 4'b1101;
	mem[2828] = 4'b1101;
	mem[2829] = 4'b1101;
	mem[2830] = 4'b1101;
	mem[2831] = 4'b1101;
	mem[2832] = 4'b1101;
	mem[2833] = 4'b1101;
	mem[2834] = 4'b1101;
	mem[2835] = 4'b1101;
	mem[2836] = 4'b0111;
	mem[2837] = 4'b0101;
	mem[2838] = 4'b0101;
	mem[2839] = 4'b0101;
	mem[2840] = 4'b0101;
	mem[2841] = 4'b0101;
	mem[2842] = 4'b0101;
	mem[2843] = 4'b0101;
	mem[2844] = 4'b0101;
	mem[2845] = 4'b0101;
	mem[2846] = 4'b0101;
	mem[2847] = 4'b0101;
	mem[2848] = 4'b0101;
	mem[2849] = 4'b0101;
	mem[2850] = 4'b0101;
	mem[2851] = 4'b0101;
	mem[2852] = 4'b0101;
	mem[2853] = 4'b1101;
	mem[2854] = 4'b1111;
	mem[2855] = 4'b1111;
	mem[2856] = 4'b1111;
	mem[2857] = 4'b1111;
	mem[2858] = 4'b1111;
	mem[2859] = 4'b1111;
	mem[2860] = 4'b1111;
	mem[2861] = 4'b1111;
	mem[2862] = 4'b1111;
	mem[2863] = 4'b1111;
	mem[2864] = 4'b1111;
	mem[2865] = 4'b1110;
	mem[2866] = 4'b1101;
	mem[2867] = 4'b1110;
	mem[2868] = 4'b1110;
	mem[2869] = 4'b1101;
	mem[2870] = 4'b1000;
	mem[2871] = 4'b0110;
	mem[2872] = 4'b0110;
	mem[2873] = 4'b0110;
	mem[2874] = 4'b0110;
	mem[2875] = 4'b0101;
	mem[2876] = 4'b0101;
	mem[2877] = 4'b0110;
	mem[2878] = 4'b0110;
	mem[2879] = 4'b0110;
	mem[2880] = 4'b0110;
	mem[2881] = 4'b0110;
	mem[2882] = 4'b0110;
	mem[2883] = 4'b0110;
	mem[2884] = 4'b0110;
	mem[2885] = 4'b0110;
	mem[2886] = 4'b0110;
	mem[2887] = 4'b1101;
	mem[2888] = 4'b1111;
	mem[2889] = 4'b1111;
	mem[2890] = 4'b1111;
	mem[2891] = 4'b1111;
	mem[2892] = 4'b1111;
	mem[2893] = 4'b1111;
	mem[2894] = 4'b1111;
	mem[2895] = 4'b1111;
	mem[2896] = 4'b1111;
	mem[2897] = 4'b1111;
	mem[2898] = 4'b1111;
	mem[2899] = 4'b1111;
	mem[2900] = 4'b1111;
	mem[2901] = 4'b1111;
	mem[2902] = 4'b1111;
	mem[2903] = 4'b1111;
	mem[2904] = 4'b1001;
	mem[2905] = 4'b0110;
	mem[2906] = 4'b0110;
	mem[2907] = 4'b0110;
	mem[2908] = 4'b0110;
	mem[2909] = 4'b0110;
	mem[2910] = 4'b0110;
	mem[2911] = 4'b0110;
	mem[2912] = 4'b0110;
	mem[2913] = 4'b0110;
	mem[2914] = 4'b0110;
	mem[2915] = 4'b0110;
	mem[2916] = 4'b0110;
	mem[2917] = 4'b0110;
	mem[2918] = 4'b0111;
	mem[2919] = 4'b0111;
	mem[2920] = 4'b0111;
	mem[2921] = 4'b1100;
	mem[2922] = 4'b1111;
	mem[2923] = 4'b1111;
	mem[2924] = 4'b1101;
	mem[2925] = 4'b1101;
	mem[2926] = 4'b1101;
	mem[2927] = 4'b1101;
	mem[2928] = 4'b1101;
	mem[2929] = 4'b1101;
	mem[2930] = 4'b1101;
	mem[2931] = 4'b1101;
	mem[2932] = 4'b1101;
	mem[2933] = 4'b1101;
	mem[2934] = 4'b1111;
	mem[2935] = 4'b1111;
	mem[2936] = 4'b1111;
	mem[2937] = 4'b1111;
	mem[2938] = 4'b0011;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b0111;
	mem[2948] = 4'b1100;
	mem[2949] = 4'b1101;
	mem[2950] = 4'b1101;
	mem[2951] = 4'b1101;
	mem[2952] = 4'b1101;
	mem[2953] = 4'b1101;
	mem[2954] = 4'b1101;
	mem[2955] = 4'b1101;
	mem[2956] = 4'b1101;
	mem[2957] = 4'b1101;
	mem[2958] = 4'b1101;
	mem[2959] = 4'b1101;
	mem[2960] = 4'b1101;
	mem[2961] = 4'b1101;
	mem[2962] = 4'b1101;
	mem[2963] = 4'b1101;
	mem[2964] = 4'b0111;
	mem[2965] = 4'b0101;
	mem[2966] = 4'b0101;
	mem[2967] = 4'b0101;
	mem[2968] = 4'b0101;
	mem[2969] = 4'b0101;
	mem[2970] = 4'b0101;
	mem[2971] = 4'b0101;
	mem[2972] = 4'b0101;
	mem[2973] = 4'b0101;
	mem[2974] = 4'b0101;
	mem[2975] = 4'b0101;
	mem[2976] = 4'b0101;
	mem[2977] = 4'b0101;
	mem[2978] = 4'b0101;
	mem[2979] = 4'b0101;
	mem[2980] = 4'b0101;
	mem[2981] = 4'b1101;
	mem[2982] = 4'b1111;
	mem[2983] = 4'b1111;
	mem[2984] = 4'b1111;
	mem[2985] = 4'b1111;
	mem[2986] = 4'b1111;
	mem[2987] = 4'b1111;
	mem[2988] = 4'b1111;
	mem[2989] = 4'b1111;
	mem[2990] = 4'b1111;
	mem[2991] = 4'b1111;
	mem[2992] = 4'b1111;
	mem[2993] = 4'b1101;
	mem[2994] = 4'b1110;
	mem[2995] = 4'b1111;
	mem[2996] = 4'b1111;
	mem[2997] = 4'b1101;
	mem[2998] = 4'b1000;
	mem[2999] = 4'b0101;
	mem[3000] = 4'b0110;
	mem[3001] = 4'b0110;
	mem[3002] = 4'b0110;
	mem[3003] = 4'b0110;
	mem[3004] = 4'b0110;
	mem[3005] = 4'b0110;
	mem[3006] = 4'b0110;
	mem[3007] = 4'b0110;
	mem[3008] = 4'b0110;
	mem[3009] = 4'b0110;
	mem[3010] = 4'b0110;
	mem[3011] = 4'b0110;
	mem[3012] = 4'b0110;
	mem[3013] = 4'b0110;
	mem[3014] = 4'b0110;
	mem[3015] = 4'b1101;
	mem[3016] = 4'b1111;
	mem[3017] = 4'b1111;
	mem[3018] = 4'b1111;
	mem[3019] = 4'b1111;
	mem[3020] = 4'b1111;
	mem[3021] = 4'b1111;
	mem[3022] = 4'b1111;
	mem[3023] = 4'b1111;
	mem[3024] = 4'b1111;
	mem[3025] = 4'b1111;
	mem[3026] = 4'b1111;
	mem[3027] = 4'b1111;
	mem[3028] = 4'b1111;
	mem[3029] = 4'b1111;
	mem[3030] = 4'b1111;
	mem[3031] = 4'b1111;
	mem[3032] = 4'b1001;
	mem[3033] = 4'b0110;
	mem[3034] = 4'b0110;
	mem[3035] = 4'b0110;
	mem[3036] = 4'b0110;
	mem[3037] = 4'b0110;
	mem[3038] = 4'b0110;
	mem[3039] = 4'b0110;
	mem[3040] = 4'b0110;
	mem[3041] = 4'b0110;
	mem[3042] = 4'b0110;
	mem[3043] = 4'b0110;
	mem[3044] = 4'b0110;
	mem[3045] = 4'b0110;
	mem[3046] = 4'b0110;
	mem[3047] = 4'b0110;
	mem[3048] = 4'b0111;
	mem[3049] = 4'b1100;
	mem[3050] = 4'b1111;
	mem[3051] = 4'b1111;
	mem[3052] = 4'b1111;
	mem[3053] = 4'b1110;
	mem[3054] = 4'b1101;
	mem[3055] = 4'b1101;
	mem[3056] = 4'b1101;
	mem[3057] = 4'b1101;
	mem[3058] = 4'b1101;
	mem[3059] = 4'b1101;
	mem[3060] = 4'b1101;
	mem[3061] = 4'b1111;
	mem[3062] = 4'b1111;
	mem[3063] = 4'b1111;
	mem[3064] = 4'b1111;
	mem[3065] = 4'b1111;
	mem[3066] = 4'b0011;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b0111;
	mem[3076] = 4'b1100;
	mem[3077] = 4'b1101;
	mem[3078] = 4'b1101;
	mem[3079] = 4'b1101;
	mem[3080] = 4'b1101;
	mem[3081] = 4'b1101;
	mem[3082] = 4'b1101;
	mem[3083] = 4'b1101;
	mem[3084] = 4'b1101;
	mem[3085] = 4'b1101;
	mem[3086] = 4'b1101;
	mem[3087] = 4'b1101;
	mem[3088] = 4'b1101;
	mem[3089] = 4'b1101;
	mem[3090] = 4'b1101;
	mem[3091] = 4'b1101;
	mem[3092] = 4'b0111;
	mem[3093] = 4'b0101;
	mem[3094] = 4'b0101;
	mem[3095] = 4'b0101;
	mem[3096] = 4'b0101;
	mem[3097] = 4'b0101;
	mem[3098] = 4'b0101;
	mem[3099] = 4'b0101;
	mem[3100] = 4'b0101;
	mem[3101] = 4'b0101;
	mem[3102] = 4'b0101;
	mem[3103] = 4'b0101;
	mem[3104] = 4'b0101;
	mem[3105] = 4'b0101;
	mem[3106] = 4'b0101;
	mem[3107] = 4'b0101;
	mem[3108] = 4'b0101;
	mem[3109] = 4'b1101;
	mem[3110] = 4'b1111;
	mem[3111] = 4'b1111;
	mem[3112] = 4'b1111;
	mem[3113] = 4'b1111;
	mem[3114] = 4'b1111;
	mem[3115] = 4'b1111;
	mem[3116] = 4'b1111;
	mem[3117] = 4'b1111;
	mem[3118] = 4'b1111;
	mem[3119] = 4'b1111;
	mem[3120] = 4'b1110;
	mem[3121] = 4'b1101;
	mem[3122] = 4'b1111;
	mem[3123] = 4'b1111;
	mem[3124] = 4'b1110;
	mem[3125] = 4'b1110;
	mem[3126] = 4'b1001;
	mem[3127] = 4'b0101;
	mem[3128] = 4'b0101;
	mem[3129] = 4'b0110;
	mem[3130] = 4'b0110;
	mem[3131] = 4'b0110;
	mem[3132] = 4'b0110;
	mem[3133] = 4'b0110;
	mem[3134] = 4'b0110;
	mem[3135] = 4'b0110;
	mem[3136] = 4'b0110;
	mem[3137] = 4'b0110;
	mem[3138] = 4'b0110;
	mem[3139] = 4'b0110;
	mem[3140] = 4'b0110;
	mem[3141] = 4'b0110;
	mem[3142] = 4'b0110;
	mem[3143] = 4'b1101;
	mem[3144] = 4'b1111;
	mem[3145] = 4'b1111;
	mem[3146] = 4'b1111;
	mem[3147] = 4'b1111;
	mem[3148] = 4'b1111;
	mem[3149] = 4'b1111;
	mem[3150] = 4'b1111;
	mem[3151] = 4'b1111;
	mem[3152] = 4'b1111;
	mem[3153] = 4'b1111;
	mem[3154] = 4'b1111;
	mem[3155] = 4'b1111;
	mem[3156] = 4'b1111;
	mem[3157] = 4'b1111;
	mem[3158] = 4'b1111;
	mem[3159] = 4'b1111;
	mem[3160] = 4'b1001;
	mem[3161] = 4'b0110;
	mem[3162] = 4'b0110;
	mem[3163] = 4'b0110;
	mem[3164] = 4'b0110;
	mem[3165] = 4'b0110;
	mem[3166] = 4'b0110;
	mem[3167] = 4'b0110;
	mem[3168] = 4'b0110;
	mem[3169] = 4'b0110;
	mem[3170] = 4'b0110;
	mem[3171] = 4'b0110;
	mem[3172] = 4'b0110;
	mem[3173] = 4'b0110;
	mem[3174] = 4'b0110;
	mem[3175] = 4'b0110;
	mem[3176] = 4'b0110;
	mem[3177] = 4'b1100;
	mem[3178] = 4'b1111;
	mem[3179] = 4'b1111;
	mem[3180] = 4'b1111;
	mem[3181] = 4'b1111;
	mem[3182] = 4'b1111;
	mem[3183] = 4'b1110;
	mem[3184] = 4'b1101;
	mem[3185] = 4'b1101;
	mem[3186] = 4'b1101;
	mem[3187] = 4'b1110;
	mem[3188] = 4'b1111;
	mem[3189] = 4'b1111;
	mem[3190] = 4'b1111;
	mem[3191] = 4'b1111;
	mem[3192] = 4'b1111;
	mem[3193] = 4'b1111;
	mem[3194] = 4'b0011;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b0111;
	mem[3204] = 4'b1100;
	mem[3205] = 4'b1101;
	mem[3206] = 4'b1101;
	mem[3207] = 4'b1101;
	mem[3208] = 4'b1101;
	mem[3209] = 4'b1101;
	mem[3210] = 4'b1101;
	mem[3211] = 4'b1101;
	mem[3212] = 4'b1101;
	mem[3213] = 4'b1101;
	mem[3214] = 4'b1101;
	mem[3215] = 4'b1101;
	mem[3216] = 4'b1101;
	mem[3217] = 4'b1101;
	mem[3218] = 4'b1101;
	mem[3219] = 4'b1101;
	mem[3220] = 4'b0111;
	mem[3221] = 4'b0101;
	mem[3222] = 4'b0101;
	mem[3223] = 4'b0101;
	mem[3224] = 4'b0101;
	mem[3225] = 4'b0101;
	mem[3226] = 4'b0101;
	mem[3227] = 4'b0101;
	mem[3228] = 4'b0101;
	mem[3229] = 4'b0101;
	mem[3230] = 4'b0101;
	mem[3231] = 4'b0101;
	mem[3232] = 4'b0101;
	mem[3233] = 4'b0101;
	mem[3234] = 4'b0101;
	mem[3235] = 4'b0101;
	mem[3236] = 4'b0101;
	mem[3237] = 4'b1101;
	mem[3238] = 4'b1111;
	mem[3239] = 4'b1111;
	mem[3240] = 4'b1111;
	mem[3241] = 4'b1111;
	mem[3242] = 4'b1111;
	mem[3243] = 4'b1111;
	mem[3244] = 4'b1111;
	mem[3245] = 4'b1111;
	mem[3246] = 4'b1111;
	mem[3247] = 4'b1111;
	mem[3248] = 4'b1111;
	mem[3249] = 4'b1110;
	mem[3250] = 4'b1111;
	mem[3251] = 4'b1111;
	mem[3252] = 4'b1101;
	mem[3253] = 4'b1111;
	mem[3254] = 4'b1010;
	mem[3255] = 4'b0101;
	mem[3256] = 4'b0101;
	mem[3257] = 4'b0101;
	mem[3258] = 4'b0110;
	mem[3259] = 4'b0110;
	mem[3260] = 4'b0110;
	mem[3261] = 4'b0110;
	mem[3262] = 4'b0110;
	mem[3263] = 4'b0110;
	mem[3264] = 4'b0110;
	mem[3265] = 4'b0110;
	mem[3266] = 4'b0110;
	mem[3267] = 4'b0110;
	mem[3268] = 4'b0110;
	mem[3269] = 4'b0110;
	mem[3270] = 4'b0110;
	mem[3271] = 4'b1101;
	mem[3272] = 4'b1111;
	mem[3273] = 4'b1111;
	mem[3274] = 4'b1111;
	mem[3275] = 4'b1111;
	mem[3276] = 4'b1111;
	mem[3277] = 4'b1111;
	mem[3278] = 4'b1111;
	mem[3279] = 4'b1111;
	mem[3280] = 4'b1111;
	mem[3281] = 4'b1111;
	mem[3282] = 4'b1111;
	mem[3283] = 4'b1111;
	mem[3284] = 4'b1111;
	mem[3285] = 4'b1111;
	mem[3286] = 4'b1111;
	mem[3287] = 4'b1111;
	mem[3288] = 4'b1001;
	mem[3289] = 4'b0110;
	mem[3290] = 4'b0110;
	mem[3291] = 4'b0110;
	mem[3292] = 4'b0110;
	mem[3293] = 4'b0110;
	mem[3294] = 4'b0110;
	mem[3295] = 4'b0110;
	mem[3296] = 4'b0110;
	mem[3297] = 4'b0110;
	mem[3298] = 4'b0111;
	mem[3299] = 4'b0111;
	mem[3300] = 4'b0110;
	mem[3301] = 4'b0110;
	mem[3302] = 4'b0110;
	mem[3303] = 4'b0110;
	mem[3304] = 4'b0110;
	mem[3305] = 4'b1011;
	mem[3306] = 4'b1111;
	mem[3307] = 4'b1111;
	mem[3308] = 4'b1111;
	mem[3309] = 4'b1111;
	mem[3310] = 4'b1111;
	mem[3311] = 4'b1111;
	mem[3312] = 4'b1111;
	mem[3313] = 4'b1111;
	mem[3314] = 4'b1111;
	mem[3315] = 4'b1111;
	mem[3316] = 4'b1111;
	mem[3317] = 4'b1111;
	mem[3318] = 4'b1111;
	mem[3319] = 4'b1111;
	mem[3320] = 4'b1111;
	mem[3321] = 4'b1111;
	mem[3322] = 4'b0011;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b0111;
	mem[3332] = 4'b1100;
	mem[3333] = 4'b1101;
	mem[3334] = 4'b1101;
	mem[3335] = 4'b1101;
	mem[3336] = 4'b1101;
	mem[3337] = 4'b1101;
	mem[3338] = 4'b1101;
	mem[3339] = 4'b1101;
	mem[3340] = 4'b1101;
	mem[3341] = 4'b1101;
	mem[3342] = 4'b1101;
	mem[3343] = 4'b1101;
	mem[3344] = 4'b1101;
	mem[3345] = 4'b1101;
	mem[3346] = 4'b1101;
	mem[3347] = 4'b1101;
	mem[3348] = 4'b0111;
	mem[3349] = 4'b0101;
	mem[3350] = 4'b0101;
	mem[3351] = 4'b0101;
	mem[3352] = 4'b0101;
	mem[3353] = 4'b0101;
	mem[3354] = 4'b0101;
	mem[3355] = 4'b0101;
	mem[3356] = 4'b0101;
	mem[3357] = 4'b0101;
	mem[3358] = 4'b0101;
	mem[3359] = 4'b0101;
	mem[3360] = 4'b0101;
	mem[3361] = 4'b0101;
	mem[3362] = 4'b0101;
	mem[3363] = 4'b0101;
	mem[3364] = 4'b0101;
	mem[3365] = 4'b1101;
	mem[3366] = 4'b1111;
	mem[3367] = 4'b1111;
	mem[3368] = 4'b1111;
	mem[3369] = 4'b1111;
	mem[3370] = 4'b1111;
	mem[3371] = 4'b1111;
	mem[3372] = 4'b1111;
	mem[3373] = 4'b1111;
	mem[3374] = 4'b1111;
	mem[3375] = 4'b1111;
	mem[3376] = 4'b1111;
	mem[3377] = 4'b1111;
	mem[3378] = 4'b1111;
	mem[3379] = 4'b1110;
	mem[3380] = 4'b1110;
	mem[3381] = 4'b1111;
	mem[3382] = 4'b1001;
	mem[3383] = 4'b0101;
	mem[3384] = 4'b0101;
	mem[3385] = 4'b0110;
	mem[3386] = 4'b0111;
	mem[3387] = 4'b0110;
	mem[3388] = 4'b0110;
	mem[3389] = 4'b0110;
	mem[3390] = 4'b0110;
	mem[3391] = 4'b0110;
	mem[3392] = 4'b0110;
	mem[3393] = 4'b0110;
	mem[3394] = 4'b0110;
	mem[3395] = 4'b0110;
	mem[3396] = 4'b0110;
	mem[3397] = 4'b0110;
	mem[3398] = 4'b0110;
	mem[3399] = 4'b1101;
	mem[3400] = 4'b1111;
	mem[3401] = 4'b1111;
	mem[3402] = 4'b1111;
	mem[3403] = 4'b1111;
	mem[3404] = 4'b1111;
	mem[3405] = 4'b1111;
	mem[3406] = 4'b1111;
	mem[3407] = 4'b1111;
	mem[3408] = 4'b1111;
	mem[3409] = 4'b1111;
	mem[3410] = 4'b1111;
	mem[3411] = 4'b1111;
	mem[3412] = 4'b1111;
	mem[3413] = 4'b1111;
	mem[3414] = 4'b1111;
	mem[3415] = 4'b1111;
	mem[3416] = 4'b1001;
	mem[3417] = 4'b0110;
	mem[3418] = 4'b0110;
	mem[3419] = 4'b0110;
	mem[3420] = 4'b0110;
	mem[3421] = 4'b0110;
	mem[3422] = 4'b0110;
	mem[3423] = 4'b0110;
	mem[3424] = 4'b0110;
	mem[3425] = 4'b0111;
	mem[3426] = 4'b0111;
	mem[3427] = 4'b0111;
	mem[3428] = 4'b0111;
	mem[3429] = 4'b0110;
	mem[3430] = 4'b0110;
	mem[3431] = 4'b0110;
	mem[3432] = 4'b0110;
	mem[3433] = 4'b1011;
	mem[3434] = 4'b1110;
	mem[3435] = 4'b1111;
	mem[3436] = 4'b1111;
	mem[3437] = 4'b1111;
	mem[3438] = 4'b1111;
	mem[3439] = 4'b1111;
	mem[3440] = 4'b1111;
	mem[3441] = 4'b1111;
	mem[3442] = 4'b1111;
	mem[3443] = 4'b1111;
	mem[3444] = 4'b1111;
	mem[3445] = 4'b1111;
	mem[3446] = 4'b1111;
	mem[3447] = 4'b1111;
	mem[3448] = 4'b1111;
	mem[3449] = 4'b1111;
	mem[3450] = 4'b0011;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b0111;
	mem[3460] = 4'b1100;
	mem[3461] = 4'b1101;
	mem[3462] = 4'b1101;
	mem[3463] = 4'b1101;
	mem[3464] = 4'b1101;
	mem[3465] = 4'b1101;
	mem[3466] = 4'b1101;
	mem[3467] = 4'b1101;
	mem[3468] = 4'b1101;
	mem[3469] = 4'b1101;
	mem[3470] = 4'b1101;
	mem[3471] = 4'b1101;
	mem[3472] = 4'b1101;
	mem[3473] = 4'b1101;
	mem[3474] = 4'b1101;
	mem[3475] = 4'b1101;
	mem[3476] = 4'b0111;
	mem[3477] = 4'b0101;
	mem[3478] = 4'b0101;
	mem[3479] = 4'b0101;
	mem[3480] = 4'b0101;
	mem[3481] = 4'b0101;
	mem[3482] = 4'b0101;
	mem[3483] = 4'b0101;
	mem[3484] = 4'b0101;
	mem[3485] = 4'b0101;
	mem[3486] = 4'b0101;
	mem[3487] = 4'b0101;
	mem[3488] = 4'b0101;
	mem[3489] = 4'b0101;
	mem[3490] = 4'b0101;
	mem[3491] = 4'b0101;
	mem[3492] = 4'b0101;
	mem[3493] = 4'b1101;
	mem[3494] = 4'b1111;
	mem[3495] = 4'b1111;
	mem[3496] = 4'b1111;
	mem[3497] = 4'b1111;
	mem[3498] = 4'b1111;
	mem[3499] = 4'b1111;
	mem[3500] = 4'b1111;
	mem[3501] = 4'b1111;
	mem[3502] = 4'b1111;
	mem[3503] = 4'b1111;
	mem[3504] = 4'b1111;
	mem[3505] = 4'b1111;
	mem[3506] = 4'b1111;
	mem[3507] = 4'b1101;
	mem[3508] = 4'b1110;
	mem[3509] = 4'b1111;
	mem[3510] = 4'b1001;
	mem[3511] = 4'b0101;
	mem[3512] = 4'b0110;
	mem[3513] = 4'b0110;
	mem[3514] = 4'b0110;
	mem[3515] = 4'b0110;
	mem[3516] = 4'b0110;
	mem[3517] = 4'b0110;
	mem[3518] = 4'b0110;
	mem[3519] = 4'b0110;
	mem[3520] = 4'b0110;
	mem[3521] = 4'b0110;
	mem[3522] = 4'b0110;
	mem[3523] = 4'b0110;
	mem[3524] = 4'b0110;
	mem[3525] = 4'b0110;
	mem[3526] = 4'b0110;
	mem[3527] = 4'b1101;
	mem[3528] = 4'b1111;
	mem[3529] = 4'b1111;
	mem[3530] = 4'b1111;
	mem[3531] = 4'b1111;
	mem[3532] = 4'b1111;
	mem[3533] = 4'b1111;
	mem[3534] = 4'b1111;
	mem[3535] = 4'b1111;
	mem[3536] = 4'b1111;
	mem[3537] = 4'b1111;
	mem[3538] = 4'b1111;
	mem[3539] = 4'b1111;
	mem[3540] = 4'b1111;
	mem[3541] = 4'b1111;
	mem[3542] = 4'b1111;
	mem[3543] = 4'b1111;
	mem[3544] = 4'b1001;
	mem[3545] = 4'b0110;
	mem[3546] = 4'b0110;
	mem[3547] = 4'b0110;
	mem[3548] = 4'b0110;
	mem[3549] = 4'b0110;
	mem[3550] = 4'b0111;
	mem[3551] = 4'b0110;
	mem[3552] = 4'b0111;
	mem[3553] = 4'b0111;
	mem[3554] = 4'b0111;
	mem[3555] = 4'b0111;
	mem[3556] = 4'b0111;
	mem[3557] = 4'b0111;
	mem[3558] = 4'b0110;
	mem[3559] = 4'b0110;
	mem[3560] = 4'b0110;
	mem[3561] = 4'b1011;
	mem[3562] = 4'b1101;
	mem[3563] = 4'b1110;
	mem[3564] = 4'b1111;
	mem[3565] = 4'b1111;
	mem[3566] = 4'b1111;
	mem[3567] = 4'b1111;
	mem[3568] = 4'b1111;
	mem[3569] = 4'b1111;
	mem[3570] = 4'b1111;
	mem[3571] = 4'b1111;
	mem[3572] = 4'b1111;
	mem[3573] = 4'b1111;
	mem[3574] = 4'b1111;
	mem[3575] = 4'b1111;
	mem[3576] = 4'b1111;
	mem[3577] = 4'b1111;
	mem[3578] = 4'b0011;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b0111;
	mem[3588] = 4'b1100;
	mem[3589] = 4'b1101;
	mem[3590] = 4'b1101;
	mem[3591] = 4'b1101;
	mem[3592] = 4'b1101;
	mem[3593] = 4'b1101;
	mem[3594] = 4'b1101;
	mem[3595] = 4'b1101;
	mem[3596] = 4'b1101;
	mem[3597] = 4'b1101;
	mem[3598] = 4'b1101;
	mem[3599] = 4'b1101;
	mem[3600] = 4'b1101;
	mem[3601] = 4'b1101;
	mem[3602] = 4'b1101;
	mem[3603] = 4'b1101;
	mem[3604] = 4'b0111;
	mem[3605] = 4'b0101;
	mem[3606] = 4'b0101;
	mem[3607] = 4'b0101;
	mem[3608] = 4'b0101;
	mem[3609] = 4'b0101;
	mem[3610] = 4'b0101;
	mem[3611] = 4'b0101;
	mem[3612] = 4'b0101;
	mem[3613] = 4'b0101;
	mem[3614] = 4'b0101;
	mem[3615] = 4'b0101;
	mem[3616] = 4'b0101;
	mem[3617] = 4'b0101;
	mem[3618] = 4'b0101;
	mem[3619] = 4'b0101;
	mem[3620] = 4'b0101;
	mem[3621] = 4'b1101;
	mem[3622] = 4'b1111;
	mem[3623] = 4'b1101;
	mem[3624] = 4'b1110;
	mem[3625] = 4'b1111;
	mem[3626] = 4'b1111;
	mem[3627] = 4'b1111;
	mem[3628] = 4'b1111;
	mem[3629] = 4'b1111;
	mem[3630] = 4'b1111;
	mem[3631] = 4'b1111;
	mem[3632] = 4'b1111;
	mem[3633] = 4'b1111;
	mem[3634] = 4'b1111;
	mem[3635] = 4'b1101;
	mem[3636] = 4'b1101;
	mem[3637] = 4'b1101;
	mem[3638] = 4'b1000;
	mem[3639] = 4'b0110;
	mem[3640] = 4'b0111;
	mem[3641] = 4'b0110;
	mem[3642] = 4'b0110;
	mem[3643] = 4'b0110;
	mem[3644] = 4'b0110;
	mem[3645] = 4'b0110;
	mem[3646] = 4'b0110;
	mem[3647] = 4'b0110;
	mem[3648] = 4'b0110;
	mem[3649] = 4'b0110;
	mem[3650] = 4'b0110;
	mem[3651] = 4'b0110;
	mem[3652] = 4'b0110;
	mem[3653] = 4'b0110;
	mem[3654] = 4'b0110;
	mem[3655] = 4'b1101;
	mem[3656] = 4'b1111;
	mem[3657] = 4'b1111;
	mem[3658] = 4'b1111;
	mem[3659] = 4'b1111;
	mem[3660] = 4'b1111;
	mem[3661] = 4'b1111;
	mem[3662] = 4'b1111;
	mem[3663] = 4'b1111;
	mem[3664] = 4'b1111;
	mem[3665] = 4'b1111;
	mem[3666] = 4'b1111;
	mem[3667] = 4'b1111;
	mem[3668] = 4'b1111;
	mem[3669] = 4'b1111;
	mem[3670] = 4'b1111;
	mem[3671] = 4'b1111;
	mem[3672] = 4'b1001;
	mem[3673] = 4'b0110;
	mem[3674] = 4'b0110;
	mem[3675] = 4'b0110;
	mem[3676] = 4'b0110;
	mem[3677] = 4'b0110;
	mem[3678] = 4'b0110;
	mem[3679] = 4'b0110;
	mem[3680] = 4'b0111;
	mem[3681] = 4'b0111;
	mem[3682] = 4'b0111;
	mem[3683] = 4'b0111;
	mem[3684] = 4'b0111;
	mem[3685] = 4'b0111;
	mem[3686] = 4'b0111;
	mem[3687] = 4'b0111;
	mem[3688] = 4'b0110;
	mem[3689] = 4'b1011;
	mem[3690] = 4'b1101;
	mem[3691] = 4'b1101;
	mem[3692] = 4'b1110;
	mem[3693] = 4'b1111;
	mem[3694] = 4'b1111;
	mem[3695] = 4'b1111;
	mem[3696] = 4'b1111;
	mem[3697] = 4'b1111;
	mem[3698] = 4'b1111;
	mem[3699] = 4'b1111;
	mem[3700] = 4'b1111;
	mem[3701] = 4'b1111;
	mem[3702] = 4'b1111;
	mem[3703] = 4'b1111;
	mem[3704] = 4'b1111;
	mem[3705] = 4'b1111;
	mem[3706] = 4'b0011;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b0111;
	mem[3716] = 4'b1100;
	mem[3717] = 4'b1101;
	mem[3718] = 4'b1101;
	mem[3719] = 4'b1101;
	mem[3720] = 4'b1101;
	mem[3721] = 4'b1101;
	mem[3722] = 4'b1101;
	mem[3723] = 4'b1101;
	mem[3724] = 4'b1101;
	mem[3725] = 4'b1101;
	mem[3726] = 4'b1101;
	mem[3727] = 4'b1101;
	mem[3728] = 4'b1101;
	mem[3729] = 4'b1101;
	mem[3730] = 4'b1101;
	mem[3731] = 4'b1101;
	mem[3732] = 4'b0111;
	mem[3733] = 4'b0101;
	mem[3734] = 4'b0101;
	mem[3735] = 4'b0101;
	mem[3736] = 4'b0101;
	mem[3737] = 4'b0101;
	mem[3738] = 4'b0101;
	mem[3739] = 4'b0101;
	mem[3740] = 4'b0101;
	mem[3741] = 4'b0101;
	mem[3742] = 4'b0101;
	mem[3743] = 4'b0101;
	mem[3744] = 4'b0101;
	mem[3745] = 4'b0101;
	mem[3746] = 4'b0101;
	mem[3747] = 4'b0101;
	mem[3748] = 4'b0101;
	mem[3749] = 4'b1101;
	mem[3750] = 4'b1110;
	mem[3751] = 4'b1101;
	mem[3752] = 4'b1101;
	mem[3753] = 4'b1110;
	mem[3754] = 4'b1111;
	mem[3755] = 4'b1111;
	mem[3756] = 4'b1111;
	mem[3757] = 4'b1111;
	mem[3758] = 4'b1111;
	mem[3759] = 4'b1111;
	mem[3760] = 4'b1111;
	mem[3761] = 4'b1111;
	mem[3762] = 4'b1111;
	mem[3763] = 4'b1111;
	mem[3764] = 4'b1110;
	mem[3765] = 4'b1101;
	mem[3766] = 4'b1001;
	mem[3767] = 4'b0111;
	mem[3768] = 4'b0110;
	mem[3769] = 4'b0110;
	mem[3770] = 4'b0110;
	mem[3771] = 4'b0110;
	mem[3772] = 4'b0110;
	mem[3773] = 4'b0110;
	mem[3774] = 4'b0110;
	mem[3775] = 4'b0110;
	mem[3776] = 4'b0110;
	mem[3777] = 4'b0110;
	mem[3778] = 4'b0110;
	mem[3779] = 4'b0110;
	mem[3780] = 4'b0110;
	mem[3781] = 4'b0110;
	mem[3782] = 4'b0110;
	mem[3783] = 4'b1101;
	mem[3784] = 4'b1111;
	mem[3785] = 4'b1111;
	mem[3786] = 4'b1111;
	mem[3787] = 4'b1111;
	mem[3788] = 4'b1111;
	mem[3789] = 4'b1111;
	mem[3790] = 4'b1111;
	mem[3791] = 4'b1111;
	mem[3792] = 4'b1111;
	mem[3793] = 4'b1111;
	mem[3794] = 4'b1111;
	mem[3795] = 4'b1111;
	mem[3796] = 4'b1111;
	mem[3797] = 4'b1111;
	mem[3798] = 4'b1111;
	mem[3799] = 4'b1111;
	mem[3800] = 4'b1001;
	mem[3801] = 4'b0111;
	mem[3802] = 4'b0111;
	mem[3803] = 4'b0110;
	mem[3804] = 4'b0110;
	mem[3805] = 4'b0110;
	mem[3806] = 4'b0110;
	mem[3807] = 4'b0110;
	mem[3808] = 4'b0111;
	mem[3809] = 4'b0111;
	mem[3810] = 4'b0111;
	mem[3811] = 4'b0111;
	mem[3812] = 4'b0111;
	mem[3813] = 4'b0111;
	mem[3814] = 4'b0111;
	mem[3815] = 4'b0111;
	mem[3816] = 4'b0111;
	mem[3817] = 4'b1011;
	mem[3818] = 4'b1101;
	mem[3819] = 4'b1101;
	mem[3820] = 4'b1101;
	mem[3821] = 4'b1110;
	mem[3822] = 4'b1111;
	mem[3823] = 4'b1111;
	mem[3824] = 4'b1111;
	mem[3825] = 4'b1111;
	mem[3826] = 4'b1111;
	mem[3827] = 4'b1111;
	mem[3828] = 4'b1111;
	mem[3829] = 4'b1111;
	mem[3830] = 4'b1111;
	mem[3831] = 4'b1111;
	mem[3832] = 4'b1111;
	mem[3833] = 4'b1111;
	mem[3834] = 4'b0011;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b0111;
	mem[3844] = 4'b1100;
	mem[3845] = 4'b1101;
	mem[3846] = 4'b1101;
	mem[3847] = 4'b1101;
	mem[3848] = 4'b1101;
	mem[3849] = 4'b1101;
	mem[3850] = 4'b1101;
	mem[3851] = 4'b1101;
	mem[3852] = 4'b1101;
	mem[3853] = 4'b1101;
	mem[3854] = 4'b1101;
	mem[3855] = 4'b1101;
	mem[3856] = 4'b1101;
	mem[3857] = 4'b1101;
	mem[3858] = 4'b1101;
	mem[3859] = 4'b1101;
	mem[3860] = 4'b0111;
	mem[3861] = 4'b0101;
	mem[3862] = 4'b0101;
	mem[3863] = 4'b0101;
	mem[3864] = 4'b0101;
	mem[3865] = 4'b0101;
	mem[3866] = 4'b0101;
	mem[3867] = 4'b0101;
	mem[3868] = 4'b0101;
	mem[3869] = 4'b0101;
	mem[3870] = 4'b0101;
	mem[3871] = 4'b0101;
	mem[3872] = 4'b0101;
	mem[3873] = 4'b0101;
	mem[3874] = 4'b0101;
	mem[3875] = 4'b0101;
	mem[3876] = 4'b0101;
	mem[3877] = 4'b1101;
	mem[3878] = 4'b1111;
	mem[3879] = 4'b1110;
	mem[3880] = 4'b1101;
	mem[3881] = 4'b1101;
	mem[3882] = 4'b1110;
	mem[3883] = 4'b1111;
	mem[3884] = 4'b1111;
	mem[3885] = 4'b1111;
	mem[3886] = 4'b1111;
	mem[3887] = 4'b1111;
	mem[3888] = 4'b1111;
	mem[3889] = 4'b1111;
	mem[3890] = 4'b1111;
	mem[3891] = 4'b1111;
	mem[3892] = 4'b1111;
	mem[3893] = 4'b1111;
	mem[3894] = 4'b1010;
	mem[3895] = 4'b0110;
	mem[3896] = 4'b0110;
	mem[3897] = 4'b0110;
	mem[3898] = 4'b0110;
	mem[3899] = 4'b0110;
	mem[3900] = 4'b0110;
	mem[3901] = 4'b0110;
	mem[3902] = 4'b0110;
	mem[3903] = 4'b0110;
	mem[3904] = 4'b0110;
	mem[3905] = 4'b0110;
	mem[3906] = 4'b0110;
	mem[3907] = 4'b0110;
	mem[3908] = 4'b0110;
	mem[3909] = 4'b0110;
	mem[3910] = 4'b0110;
	mem[3911] = 4'b1101;
	mem[3912] = 4'b1111;
	mem[3913] = 4'b1111;
	mem[3914] = 4'b1111;
	mem[3915] = 4'b1111;
	mem[3916] = 4'b1111;
	mem[3917] = 4'b1111;
	mem[3918] = 4'b1111;
	mem[3919] = 4'b1111;
	mem[3920] = 4'b1111;
	mem[3921] = 4'b1111;
	mem[3922] = 4'b1111;
	mem[3923] = 4'b1111;
	mem[3924] = 4'b1111;
	mem[3925] = 4'b1111;
	mem[3926] = 4'b1111;
	mem[3927] = 4'b1111;
	mem[3928] = 4'b1001;
	mem[3929] = 4'b0111;
	mem[3930] = 4'b0111;
	mem[3931] = 4'b0111;
	mem[3932] = 4'b0110;
	mem[3933] = 4'b0110;
	mem[3934] = 4'b0110;
	mem[3935] = 4'b0110;
	mem[3936] = 4'b0110;
	mem[3937] = 4'b0111;
	mem[3938] = 4'b0111;
	mem[3939] = 4'b0111;
	mem[3940] = 4'b0111;
	mem[3941] = 4'b0111;
	mem[3942] = 4'b0111;
	mem[3943] = 4'b0111;
	mem[3944] = 4'b0111;
	mem[3945] = 4'b1011;
	mem[3946] = 4'b1101;
	mem[3947] = 4'b1101;
	mem[3948] = 4'b1101;
	mem[3949] = 4'b1101;
	mem[3950] = 4'b1111;
	mem[3951] = 4'b1111;
	mem[3952] = 4'b1111;
	mem[3953] = 4'b1111;
	mem[3954] = 4'b1111;
	mem[3955] = 4'b1111;
	mem[3956] = 4'b1111;
	mem[3957] = 4'b1111;
	mem[3958] = 4'b1111;
	mem[3959] = 4'b1111;
	mem[3960] = 4'b1111;
	mem[3961] = 4'b1111;
	mem[3962] = 4'b0011;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b0111;
	mem[3972] = 4'b1100;
	mem[3973] = 4'b1101;
	mem[3974] = 4'b1101;
	mem[3975] = 4'b1101;
	mem[3976] = 4'b1101;
	mem[3977] = 4'b1101;
	mem[3978] = 4'b1101;
	mem[3979] = 4'b1101;
	mem[3980] = 4'b1101;
	mem[3981] = 4'b1101;
	mem[3982] = 4'b1101;
	mem[3983] = 4'b1101;
	mem[3984] = 4'b1101;
	mem[3985] = 4'b1101;
	mem[3986] = 4'b1101;
	mem[3987] = 4'b1101;
	mem[3988] = 4'b0111;
	mem[3989] = 4'b0101;
	mem[3990] = 4'b0101;
	mem[3991] = 4'b0101;
	mem[3992] = 4'b0101;
	mem[3993] = 4'b0101;
	mem[3994] = 4'b0101;
	mem[3995] = 4'b0101;
	mem[3996] = 4'b0101;
	mem[3997] = 4'b0101;
	mem[3998] = 4'b0101;
	mem[3999] = 4'b0101;
	mem[4000] = 4'b0101;
	mem[4001] = 4'b0101;
	mem[4002] = 4'b0101;
	mem[4003] = 4'b0101;
	mem[4004] = 4'b0101;
	mem[4005] = 4'b1101;
	mem[4006] = 4'b1111;
	mem[4007] = 4'b1111;
	mem[4008] = 4'b1110;
	mem[4009] = 4'b1101;
	mem[4010] = 4'b1101;
	mem[4011] = 4'b1110;
	mem[4012] = 4'b1111;
	mem[4013] = 4'b1111;
	mem[4014] = 4'b1111;
	mem[4015] = 4'b1111;
	mem[4016] = 4'b1111;
	mem[4017] = 4'b1111;
	mem[4018] = 4'b1101;
	mem[4019] = 4'b1101;
	mem[4020] = 4'b1111;
	mem[4021] = 4'b1111;
	mem[4022] = 4'b1001;
	mem[4023] = 4'b0110;
	mem[4024] = 4'b0110;
	mem[4025] = 4'b0110;
	mem[4026] = 4'b0110;
	mem[4027] = 4'b0110;
	mem[4028] = 4'b0110;
	mem[4029] = 4'b0110;
	mem[4030] = 4'b0110;
	mem[4031] = 4'b0110;
	mem[4032] = 4'b0110;
	mem[4033] = 4'b0110;
	mem[4034] = 4'b0110;
	mem[4035] = 4'b0110;
	mem[4036] = 4'b0110;
	mem[4037] = 4'b0110;
	mem[4038] = 4'b0110;
	mem[4039] = 4'b1101;
	mem[4040] = 4'b1111;
	mem[4041] = 4'b1111;
	mem[4042] = 4'b1111;
	mem[4043] = 4'b1111;
	mem[4044] = 4'b1111;
	mem[4045] = 4'b1111;
	mem[4046] = 4'b1111;
	mem[4047] = 4'b1111;
	mem[4048] = 4'b1111;
	mem[4049] = 4'b1111;
	mem[4050] = 4'b1111;
	mem[4051] = 4'b1111;
	mem[4052] = 4'b1111;
	mem[4053] = 4'b1111;
	mem[4054] = 4'b1111;
	mem[4055] = 4'b1111;
	mem[4056] = 4'b1001;
	mem[4057] = 4'b0111;
	mem[4058] = 4'b0111;
	mem[4059] = 4'b0111;
	mem[4060] = 4'b0111;
	mem[4061] = 4'b0110;
	mem[4062] = 4'b0110;
	mem[4063] = 4'b0110;
	mem[4064] = 4'b0110;
	mem[4065] = 4'b0110;
	mem[4066] = 4'b0111;
	mem[4067] = 4'b0111;
	mem[4068] = 4'b0111;
	mem[4069] = 4'b0111;
	mem[4070] = 4'b0111;
	mem[4071] = 4'b0111;
	mem[4072] = 4'b0111;
	mem[4073] = 4'b1100;
	mem[4074] = 4'b1110;
	mem[4075] = 4'b1101;
	mem[4076] = 4'b1101;
	mem[4077] = 4'b1110;
	mem[4078] = 4'b1111;
	mem[4079] = 4'b1111;
	mem[4080] = 4'b1111;
	mem[4081] = 4'b1111;
	mem[4082] = 4'b1111;
	mem[4083] = 4'b1111;
	mem[4084] = 4'b1111;
	mem[4085] = 4'b1111;
	mem[4086] = 4'b1111;
	mem[4087] = 4'b1111;
	mem[4088] = 4'b1111;
	mem[4089] = 4'b1111;
	mem[4090] = 4'b0011;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_1b (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0111;
	mem[4] = 4'b1100;
	mem[5] = 4'b1101;
	mem[6] = 4'b1101;
	mem[7] = 4'b1101;
	mem[8] = 4'b1101;
	mem[9] = 4'b1101;
	mem[10] = 4'b1101;
	mem[11] = 4'b1101;
	mem[12] = 4'b1101;
	mem[13] = 4'b1101;
	mem[14] = 4'b1101;
	mem[15] = 4'b1101;
	mem[16] = 4'b1101;
	mem[17] = 4'b1101;
	mem[18] = 4'b1101;
	mem[19] = 4'b1101;
	mem[20] = 4'b0111;
	mem[21] = 4'b0101;
	mem[22] = 4'b0101;
	mem[23] = 4'b0101;
	mem[24] = 4'b0101;
	mem[25] = 4'b0101;
	mem[26] = 4'b0101;
	mem[27] = 4'b0101;
	mem[28] = 4'b0101;
	mem[29] = 4'b0101;
	mem[30] = 4'b0101;
	mem[31] = 4'b0101;
	mem[32] = 4'b0101;
	mem[33] = 4'b0101;
	mem[34] = 4'b0101;
	mem[35] = 4'b0101;
	mem[36] = 4'b0101;
	mem[37] = 4'b1101;
	mem[38] = 4'b1111;
	mem[39] = 4'b1111;
	mem[40] = 4'b1111;
	mem[41] = 4'b1110;
	mem[42] = 4'b1101;
	mem[43] = 4'b1101;
	mem[44] = 4'b1110;
	mem[45] = 4'b1111;
	mem[46] = 4'b1111;
	mem[47] = 4'b1111;
	mem[48] = 4'b1111;
	mem[49] = 4'b1101;
	mem[50] = 4'b1101;
	mem[51] = 4'b1110;
	mem[52] = 4'b1111;
	mem[53] = 4'b1111;
	mem[54] = 4'b1001;
	mem[55] = 4'b0110;
	mem[56] = 4'b0110;
	mem[57] = 4'b0110;
	mem[58] = 4'b0110;
	mem[59] = 4'b0110;
	mem[60] = 4'b0110;
	mem[61] = 4'b0110;
	mem[62] = 4'b0110;
	mem[63] = 4'b0110;
	mem[64] = 4'b0110;
	mem[65] = 4'b0110;
	mem[66] = 4'b0110;
	mem[67] = 4'b0110;
	mem[68] = 4'b0110;
	mem[69] = 4'b0110;
	mem[70] = 4'b0110;
	mem[71] = 4'b1101;
	mem[72] = 4'b1111;
	mem[73] = 4'b1111;
	mem[74] = 4'b1111;
	mem[75] = 4'b1111;
	mem[76] = 4'b1111;
	mem[77] = 4'b1111;
	mem[78] = 4'b1111;
	mem[79] = 4'b1111;
	mem[80] = 4'b1111;
	mem[81] = 4'b1111;
	mem[82] = 4'b1111;
	mem[83] = 4'b1111;
	mem[84] = 4'b1111;
	mem[85] = 4'b1111;
	mem[86] = 4'b1111;
	mem[87] = 4'b1111;
	mem[88] = 4'b1001;
	mem[89] = 4'b0111;
	mem[90] = 4'b0111;
	mem[91] = 4'b0111;
	mem[92] = 4'b0111;
	mem[93] = 4'b0111;
	mem[94] = 4'b0110;
	mem[95] = 4'b0110;
	mem[96] = 4'b0110;
	mem[97] = 4'b0110;
	mem[98] = 4'b0110;
	mem[99] = 4'b0111;
	mem[100] = 4'b0111;
	mem[101] = 4'b0111;
	mem[102] = 4'b0111;
	mem[103] = 4'b0111;
	mem[104] = 4'b0111;
	mem[105] = 4'b1100;
	mem[106] = 4'b1111;
	mem[107] = 4'b1110;
	mem[108] = 4'b1110;
	mem[109] = 4'b1111;
	mem[110] = 4'b1111;
	mem[111] = 4'b1111;
	mem[112] = 4'b1111;
	mem[113] = 4'b1111;
	mem[114] = 4'b1111;
	mem[115] = 4'b1111;
	mem[116] = 4'b1111;
	mem[117] = 4'b1111;
	mem[118] = 4'b1111;
	mem[119] = 4'b1111;
	mem[120] = 4'b1111;
	mem[121] = 4'b1111;
	mem[122] = 4'b0011;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b0111;
	mem[132] = 4'b1100;
	mem[133] = 4'b1101;
	mem[134] = 4'b1101;
	mem[135] = 4'b1101;
	mem[136] = 4'b1101;
	mem[137] = 4'b1101;
	mem[138] = 4'b1101;
	mem[139] = 4'b1101;
	mem[140] = 4'b1101;
	mem[141] = 4'b1101;
	mem[142] = 4'b1101;
	mem[143] = 4'b1101;
	mem[144] = 4'b1101;
	mem[145] = 4'b1101;
	mem[146] = 4'b1101;
	mem[147] = 4'b1101;
	mem[148] = 4'b0111;
	mem[149] = 4'b0101;
	mem[150] = 4'b0101;
	mem[151] = 4'b0101;
	mem[152] = 4'b0101;
	mem[153] = 4'b0101;
	mem[154] = 4'b0101;
	mem[155] = 4'b0101;
	mem[156] = 4'b0101;
	mem[157] = 4'b0101;
	mem[158] = 4'b0101;
	mem[159] = 4'b0101;
	mem[160] = 4'b0101;
	mem[161] = 4'b0101;
	mem[162] = 4'b0101;
	mem[163] = 4'b0101;
	mem[164] = 4'b0101;
	mem[165] = 4'b1101;
	mem[166] = 4'b1111;
	mem[167] = 4'b1111;
	mem[168] = 4'b1111;
	mem[169] = 4'b1111;
	mem[170] = 4'b1110;
	mem[171] = 4'b1101;
	mem[172] = 4'b1101;
	mem[173] = 4'b1110;
	mem[174] = 4'b1111;
	mem[175] = 4'b1111;
	mem[176] = 4'b1101;
	mem[177] = 4'b1101;
	mem[178] = 4'b1110;
	mem[179] = 4'b1111;
	mem[180] = 4'b1111;
	mem[181] = 4'b1111;
	mem[182] = 4'b1001;
	mem[183] = 4'b0110;
	mem[184] = 4'b0110;
	mem[185] = 4'b0110;
	mem[186] = 4'b0110;
	mem[187] = 4'b0110;
	mem[188] = 4'b0110;
	mem[189] = 4'b0110;
	mem[190] = 4'b0110;
	mem[191] = 4'b0110;
	mem[192] = 4'b0110;
	mem[193] = 4'b0110;
	mem[194] = 4'b0110;
	mem[195] = 4'b0110;
	mem[196] = 4'b0110;
	mem[197] = 4'b0110;
	mem[198] = 4'b0110;
	mem[199] = 4'b1101;
	mem[200] = 4'b1111;
	mem[201] = 4'b1111;
	mem[202] = 4'b1111;
	mem[203] = 4'b1111;
	mem[204] = 4'b1111;
	mem[205] = 4'b1111;
	mem[206] = 4'b1111;
	mem[207] = 4'b1111;
	mem[208] = 4'b1111;
	mem[209] = 4'b1111;
	mem[210] = 4'b1111;
	mem[211] = 4'b1111;
	mem[212] = 4'b1111;
	mem[213] = 4'b1111;
	mem[214] = 4'b1110;
	mem[215] = 4'b1110;
	mem[216] = 4'b1001;
	mem[217] = 4'b0111;
	mem[218] = 4'b0111;
	mem[219] = 4'b0111;
	mem[220] = 4'b0111;
	mem[221] = 4'b0111;
	mem[222] = 4'b0111;
	mem[223] = 4'b0110;
	mem[224] = 4'b0110;
	mem[225] = 4'b0110;
	mem[226] = 4'b0110;
	mem[227] = 4'b0110;
	mem[228] = 4'b0111;
	mem[229] = 4'b0111;
	mem[230] = 4'b0111;
	mem[231] = 4'b0111;
	mem[232] = 4'b0111;
	mem[233] = 4'b1100;
	mem[234] = 4'b1111;
	mem[235] = 4'b1111;
	mem[236] = 4'b1111;
	mem[237] = 4'b1111;
	mem[238] = 4'b1111;
	mem[239] = 4'b1111;
	mem[240] = 4'b1111;
	mem[241] = 4'b1111;
	mem[242] = 4'b1111;
	mem[243] = 4'b1111;
	mem[244] = 4'b1111;
	mem[245] = 4'b1111;
	mem[246] = 4'b1111;
	mem[247] = 4'b1111;
	mem[248] = 4'b1111;
	mem[249] = 4'b1111;
	mem[250] = 4'b0011;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0111;
	mem[260] = 4'b1100;
	mem[261] = 4'b1101;
	mem[262] = 4'b1101;
	mem[263] = 4'b1101;
	mem[264] = 4'b1101;
	mem[265] = 4'b1101;
	mem[266] = 4'b1101;
	mem[267] = 4'b1101;
	mem[268] = 4'b1101;
	mem[269] = 4'b1101;
	mem[270] = 4'b1101;
	mem[271] = 4'b1101;
	mem[272] = 4'b1101;
	mem[273] = 4'b1101;
	mem[274] = 4'b1101;
	mem[275] = 4'b1101;
	mem[276] = 4'b0111;
	mem[277] = 4'b0101;
	mem[278] = 4'b0101;
	mem[279] = 4'b0101;
	mem[280] = 4'b0101;
	mem[281] = 4'b0101;
	mem[282] = 4'b0101;
	mem[283] = 4'b0101;
	mem[284] = 4'b0101;
	mem[285] = 4'b0101;
	mem[286] = 4'b0101;
	mem[287] = 4'b0101;
	mem[288] = 4'b0101;
	mem[289] = 4'b0101;
	mem[290] = 4'b0101;
	mem[291] = 4'b0101;
	mem[292] = 4'b0101;
	mem[293] = 4'b1101;
	mem[294] = 4'b1111;
	mem[295] = 4'b1111;
	mem[296] = 4'b1111;
	mem[297] = 4'b1111;
	mem[298] = 4'b1111;
	mem[299] = 4'b1110;
	mem[300] = 4'b1101;
	mem[301] = 4'b1101;
	mem[302] = 4'b1110;
	mem[303] = 4'b1110;
	mem[304] = 4'b1101;
	mem[305] = 4'b1110;
	mem[306] = 4'b1111;
	mem[307] = 4'b1111;
	mem[308] = 4'b1111;
	mem[309] = 4'b1111;
	mem[310] = 4'b1010;
	mem[311] = 4'b0110;
	mem[312] = 4'b0110;
	mem[313] = 4'b0110;
	mem[314] = 4'b0110;
	mem[315] = 4'b0110;
	mem[316] = 4'b0110;
	mem[317] = 4'b0110;
	mem[318] = 4'b0110;
	mem[319] = 4'b0110;
	mem[320] = 4'b0110;
	mem[321] = 4'b0110;
	mem[322] = 4'b0110;
	mem[323] = 4'b0110;
	mem[324] = 4'b0110;
	mem[325] = 4'b0110;
	mem[326] = 4'b0110;
	mem[327] = 4'b1101;
	mem[328] = 4'b1111;
	mem[329] = 4'b1111;
	mem[330] = 4'b1111;
	mem[331] = 4'b1111;
	mem[332] = 4'b1111;
	mem[333] = 4'b1111;
	mem[334] = 4'b1111;
	mem[335] = 4'b1111;
	mem[336] = 4'b1111;
	mem[337] = 4'b1111;
	mem[338] = 4'b1111;
	mem[339] = 4'b1111;
	mem[340] = 4'b1110;
	mem[341] = 4'b1101;
	mem[342] = 4'b1101;
	mem[343] = 4'b1101;
	mem[344] = 4'b1000;
	mem[345] = 4'b0110;
	mem[346] = 4'b0111;
	mem[347] = 4'b0111;
	mem[348] = 4'b0111;
	mem[349] = 4'b0111;
	mem[350] = 4'b0111;
	mem[351] = 4'b0111;
	mem[352] = 4'b0110;
	mem[353] = 4'b0110;
	mem[354] = 4'b0110;
	mem[355] = 4'b0110;
	mem[356] = 4'b0110;
	mem[357] = 4'b0111;
	mem[358] = 4'b0111;
	mem[359] = 4'b0111;
	mem[360] = 4'b0111;
	mem[361] = 4'b1100;
	mem[362] = 4'b1111;
	mem[363] = 4'b1111;
	mem[364] = 4'b1111;
	mem[365] = 4'b1111;
	mem[366] = 4'b1111;
	mem[367] = 4'b1111;
	mem[368] = 4'b1111;
	mem[369] = 4'b1111;
	mem[370] = 4'b1111;
	mem[371] = 4'b1111;
	mem[372] = 4'b1111;
	mem[373] = 4'b1111;
	mem[374] = 4'b1111;
	mem[375] = 4'b1111;
	mem[376] = 4'b1111;
	mem[377] = 4'b1111;
	mem[378] = 4'b0011;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0111;
	mem[388] = 4'b1100;
	mem[389] = 4'b1101;
	mem[390] = 4'b1101;
	mem[391] = 4'b1101;
	mem[392] = 4'b1101;
	mem[393] = 4'b1101;
	mem[394] = 4'b1101;
	mem[395] = 4'b1101;
	mem[396] = 4'b1101;
	mem[397] = 4'b1101;
	mem[398] = 4'b1101;
	mem[399] = 4'b1101;
	mem[400] = 4'b1101;
	mem[401] = 4'b1101;
	mem[402] = 4'b1101;
	mem[403] = 4'b1101;
	mem[404] = 4'b0111;
	mem[405] = 4'b0101;
	mem[406] = 4'b0101;
	mem[407] = 4'b0101;
	mem[408] = 4'b0101;
	mem[409] = 4'b0101;
	mem[410] = 4'b0101;
	mem[411] = 4'b0101;
	mem[412] = 4'b0101;
	mem[413] = 4'b0101;
	mem[414] = 4'b0101;
	mem[415] = 4'b0101;
	mem[416] = 4'b0101;
	mem[417] = 4'b0101;
	mem[418] = 4'b0101;
	mem[419] = 4'b0110;
	mem[420] = 4'b0110;
	mem[421] = 4'b1101;
	mem[422] = 4'b1111;
	mem[423] = 4'b1111;
	mem[424] = 4'b1111;
	mem[425] = 4'b1110;
	mem[426] = 4'b1111;
	mem[427] = 4'b1111;
	mem[428] = 4'b1110;
	mem[429] = 4'b1101;
	mem[430] = 4'b1101;
	mem[431] = 4'b1101;
	mem[432] = 4'b1110;
	mem[433] = 4'b1111;
	mem[434] = 4'b1111;
	mem[435] = 4'b1111;
	mem[436] = 4'b1111;
	mem[437] = 4'b1111;
	mem[438] = 4'b1010;
	mem[439] = 4'b0110;
	mem[440] = 4'b0110;
	mem[441] = 4'b0110;
	mem[442] = 4'b0110;
	mem[443] = 4'b0110;
	mem[444] = 4'b0110;
	mem[445] = 4'b0110;
	mem[446] = 4'b0110;
	mem[447] = 4'b0110;
	mem[448] = 4'b0110;
	mem[449] = 4'b0110;
	mem[450] = 4'b0110;
	mem[451] = 4'b0110;
	mem[452] = 4'b0110;
	mem[453] = 4'b0110;
	mem[454] = 4'b0110;
	mem[455] = 4'b1101;
	mem[456] = 4'b1111;
	mem[457] = 4'b1111;
	mem[458] = 4'b1111;
	mem[459] = 4'b1111;
	mem[460] = 4'b1111;
	mem[461] = 4'b1111;
	mem[462] = 4'b1111;
	mem[463] = 4'b1111;
	mem[464] = 4'b1111;
	mem[465] = 4'b1111;
	mem[466] = 4'b1111;
	mem[467] = 4'b1110;
	mem[468] = 4'b1101;
	mem[469] = 4'b1101;
	mem[470] = 4'b1101;
	mem[471] = 4'b1101;
	mem[472] = 4'b1000;
	mem[473] = 4'b0110;
	mem[474] = 4'b0110;
	mem[475] = 4'b0111;
	mem[476] = 4'b0111;
	mem[477] = 4'b0111;
	mem[478] = 4'b0111;
	mem[479] = 4'b0111;
	mem[480] = 4'b0111;
	mem[481] = 4'b0110;
	mem[482] = 4'b0110;
	mem[483] = 4'b0110;
	mem[484] = 4'b0110;
	mem[485] = 4'b0110;
	mem[486] = 4'b0111;
	mem[487] = 4'b0111;
	mem[488] = 4'b0111;
	mem[489] = 4'b1100;
	mem[490] = 4'b1111;
	mem[491] = 4'b1111;
	mem[492] = 4'b1111;
	mem[493] = 4'b1111;
	mem[494] = 4'b1111;
	mem[495] = 4'b1111;
	mem[496] = 4'b1111;
	mem[497] = 4'b1111;
	mem[498] = 4'b1111;
	mem[499] = 4'b1111;
	mem[500] = 4'b1111;
	mem[501] = 4'b1111;
	mem[502] = 4'b1111;
	mem[503] = 4'b1111;
	mem[504] = 4'b1111;
	mem[505] = 4'b1111;
	mem[506] = 4'b0011;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0111;
	mem[516] = 4'b1100;
	mem[517] = 4'b1101;
	mem[518] = 4'b1101;
	mem[519] = 4'b1101;
	mem[520] = 4'b1101;
	mem[521] = 4'b1101;
	mem[522] = 4'b1101;
	mem[523] = 4'b1101;
	mem[524] = 4'b1101;
	mem[525] = 4'b1101;
	mem[526] = 4'b1101;
	mem[527] = 4'b1101;
	mem[528] = 4'b1101;
	mem[529] = 4'b1101;
	mem[530] = 4'b1101;
	mem[531] = 4'b1101;
	mem[532] = 4'b0111;
	mem[533] = 4'b0101;
	mem[534] = 4'b0101;
	mem[535] = 4'b0101;
	mem[536] = 4'b0101;
	mem[537] = 4'b0101;
	mem[538] = 4'b0101;
	mem[539] = 4'b0101;
	mem[540] = 4'b0101;
	mem[541] = 4'b0101;
	mem[542] = 4'b0101;
	mem[543] = 4'b0101;
	mem[544] = 4'b0101;
	mem[545] = 4'b0110;
	mem[546] = 4'b0110;
	mem[547] = 4'b0110;
	mem[548] = 4'b0110;
	mem[549] = 4'b1101;
	mem[550] = 4'b1111;
	mem[551] = 4'b1111;
	mem[552] = 4'b1101;
	mem[553] = 4'b1101;
	mem[554] = 4'b1110;
	mem[555] = 4'b1111;
	mem[556] = 4'b1111;
	mem[557] = 4'b1110;
	mem[558] = 4'b1101;
	mem[559] = 4'b1110;
	mem[560] = 4'b1111;
	mem[561] = 4'b1111;
	mem[562] = 4'b1111;
	mem[563] = 4'b1111;
	mem[564] = 4'b1111;
	mem[565] = 4'b1111;
	mem[566] = 4'b1010;
	mem[567] = 4'b0110;
	mem[568] = 4'b0110;
	mem[569] = 4'b0110;
	mem[570] = 4'b0110;
	mem[571] = 4'b0110;
	mem[572] = 4'b0110;
	mem[573] = 4'b0110;
	mem[574] = 4'b0110;
	mem[575] = 4'b0110;
	mem[576] = 4'b0110;
	mem[577] = 4'b0110;
	mem[578] = 4'b0110;
	mem[579] = 4'b0110;
	mem[580] = 4'b0110;
	mem[581] = 4'b0110;
	mem[582] = 4'b0110;
	mem[583] = 4'b1101;
	mem[584] = 4'b1111;
	mem[585] = 4'b1111;
	mem[586] = 4'b1111;
	mem[587] = 4'b1111;
	mem[588] = 4'b1111;
	mem[589] = 4'b1111;
	mem[590] = 4'b1111;
	mem[591] = 4'b1111;
	mem[592] = 4'b1111;
	mem[593] = 4'b1111;
	mem[594] = 4'b1110;
	mem[595] = 4'b1101;
	mem[596] = 4'b1101;
	mem[597] = 4'b1101;
	mem[598] = 4'b1101;
	mem[599] = 4'b1101;
	mem[600] = 4'b1000;
	mem[601] = 4'b0110;
	mem[602] = 4'b0110;
	mem[603] = 4'b0110;
	mem[604] = 4'b0111;
	mem[605] = 4'b0111;
	mem[606] = 4'b0111;
	mem[607] = 4'b0111;
	mem[608] = 4'b0111;
	mem[609] = 4'b0111;
	mem[610] = 4'b0110;
	mem[611] = 4'b0110;
	mem[612] = 4'b0110;
	mem[613] = 4'b0110;
	mem[614] = 4'b0111;
	mem[615] = 4'b0111;
	mem[616] = 4'b0111;
	mem[617] = 4'b1100;
	mem[618] = 4'b1111;
	mem[619] = 4'b1111;
	mem[620] = 4'b1111;
	mem[621] = 4'b1111;
	mem[622] = 4'b1111;
	mem[623] = 4'b1111;
	mem[624] = 4'b1111;
	mem[625] = 4'b1111;
	mem[626] = 4'b1111;
	mem[627] = 4'b1111;
	mem[628] = 4'b1111;
	mem[629] = 4'b1111;
	mem[630] = 4'b1111;
	mem[631] = 4'b1111;
	mem[632] = 4'b1111;
	mem[633] = 4'b1111;
	mem[634] = 4'b0011;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0111;
	mem[644] = 4'b1100;
	mem[645] = 4'b1101;
	mem[646] = 4'b1101;
	mem[647] = 4'b1101;
	mem[648] = 4'b1101;
	mem[649] = 4'b1101;
	mem[650] = 4'b1101;
	mem[651] = 4'b1101;
	mem[652] = 4'b1101;
	mem[653] = 4'b1101;
	mem[654] = 4'b1101;
	mem[655] = 4'b1101;
	mem[656] = 4'b1101;
	mem[657] = 4'b1101;
	mem[658] = 4'b1101;
	mem[659] = 4'b1101;
	mem[660] = 4'b0111;
	mem[661] = 4'b0101;
	mem[662] = 4'b0101;
	mem[663] = 4'b0101;
	mem[664] = 4'b0101;
	mem[665] = 4'b0101;
	mem[666] = 4'b0101;
	mem[667] = 4'b0101;
	mem[668] = 4'b0101;
	mem[669] = 4'b0101;
	mem[670] = 4'b0101;
	mem[671] = 4'b0110;
	mem[672] = 4'b0110;
	mem[673] = 4'b0110;
	mem[674] = 4'b0110;
	mem[675] = 4'b0110;
	mem[676] = 4'b0110;
	mem[677] = 4'b1101;
	mem[678] = 4'b1111;
	mem[679] = 4'b1101;
	mem[680] = 4'b1101;
	mem[681] = 4'b1110;
	mem[682] = 4'b1111;
	mem[683] = 4'b1111;
	mem[684] = 4'b1111;
	mem[685] = 4'b1111;
	mem[686] = 4'b1111;
	mem[687] = 4'b1111;
	mem[688] = 4'b1111;
	mem[689] = 4'b1111;
	mem[690] = 4'b1111;
	mem[691] = 4'b1111;
	mem[692] = 4'b1111;
	mem[693] = 4'b1111;
	mem[694] = 4'b1010;
	mem[695] = 4'b0110;
	mem[696] = 4'b0110;
	mem[697] = 4'b0110;
	mem[698] = 4'b0110;
	mem[699] = 4'b0110;
	mem[700] = 4'b0110;
	mem[701] = 4'b0110;
	mem[702] = 4'b0110;
	mem[703] = 4'b0110;
	mem[704] = 4'b0110;
	mem[705] = 4'b0110;
	mem[706] = 4'b0110;
	mem[707] = 4'b0110;
	mem[708] = 4'b0110;
	mem[709] = 4'b0110;
	mem[710] = 4'b0110;
	mem[711] = 4'b1101;
	mem[712] = 4'b1111;
	mem[713] = 4'b1111;
	mem[714] = 4'b1111;
	mem[715] = 4'b1111;
	mem[716] = 4'b1111;
	mem[717] = 4'b1111;
	mem[718] = 4'b1111;
	mem[719] = 4'b1111;
	mem[720] = 4'b1111;
	mem[721] = 4'b1110;
	mem[722] = 4'b1101;
	mem[723] = 4'b1101;
	mem[724] = 4'b1101;
	mem[725] = 4'b1110;
	mem[726] = 4'b1111;
	mem[727] = 4'b1111;
	mem[728] = 4'b1000;
	mem[729] = 4'b0110;
	mem[730] = 4'b0110;
	mem[731] = 4'b0110;
	mem[732] = 4'b0110;
	mem[733] = 4'b0111;
	mem[734] = 4'b0111;
	mem[735] = 4'b0111;
	mem[736] = 4'b0111;
	mem[737] = 4'b0111;
	mem[738] = 4'b0111;
	mem[739] = 4'b0110;
	mem[740] = 4'b0110;
	mem[741] = 4'b0110;
	mem[742] = 4'b0110;
	mem[743] = 4'b0111;
	mem[744] = 4'b0111;
	mem[745] = 4'b1100;
	mem[746] = 4'b1111;
	mem[747] = 4'b1111;
	mem[748] = 4'b1111;
	mem[749] = 4'b1111;
	mem[750] = 4'b1111;
	mem[751] = 4'b1111;
	mem[752] = 4'b1111;
	mem[753] = 4'b1111;
	mem[754] = 4'b1111;
	mem[755] = 4'b1111;
	mem[756] = 4'b1111;
	mem[757] = 4'b1111;
	mem[758] = 4'b1111;
	mem[759] = 4'b1111;
	mem[760] = 4'b1111;
	mem[761] = 4'b1111;
	mem[762] = 4'b0011;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0111;
	mem[772] = 4'b1100;
	mem[773] = 4'b1101;
	mem[774] = 4'b1101;
	mem[775] = 4'b1101;
	mem[776] = 4'b1101;
	mem[777] = 4'b1101;
	mem[778] = 4'b1101;
	mem[779] = 4'b1101;
	mem[780] = 4'b1101;
	mem[781] = 4'b1101;
	mem[782] = 4'b1101;
	mem[783] = 4'b1101;
	mem[784] = 4'b1101;
	mem[785] = 4'b1101;
	mem[786] = 4'b1101;
	mem[787] = 4'b1101;
	mem[788] = 4'b0111;
	mem[789] = 4'b0101;
	mem[790] = 4'b0101;
	mem[791] = 4'b0101;
	mem[792] = 4'b0101;
	mem[793] = 4'b0101;
	mem[794] = 4'b0101;
	mem[795] = 4'b0101;
	mem[796] = 4'b0101;
	mem[797] = 4'b0110;
	mem[798] = 4'b0110;
	mem[799] = 4'b0110;
	mem[800] = 4'b0101;
	mem[801] = 4'b0101;
	mem[802] = 4'b0101;
	mem[803] = 4'b0101;
	mem[804] = 4'b0110;
	mem[805] = 4'b1101;
	mem[806] = 4'b1111;
	mem[807] = 4'b1101;
	mem[808] = 4'b1110;
	mem[809] = 4'b1111;
	mem[810] = 4'b1111;
	mem[811] = 4'b1111;
	mem[812] = 4'b1111;
	mem[813] = 4'b1111;
	mem[814] = 4'b1111;
	mem[815] = 4'b1111;
	mem[816] = 4'b1111;
	mem[817] = 4'b1111;
	mem[818] = 4'b1111;
	mem[819] = 4'b1111;
	mem[820] = 4'b1111;
	mem[821] = 4'b1111;
	mem[822] = 4'b1010;
	mem[823] = 4'b0110;
	mem[824] = 4'b0110;
	mem[825] = 4'b0110;
	mem[826] = 4'b0110;
	mem[827] = 4'b0110;
	mem[828] = 4'b0110;
	mem[829] = 4'b0110;
	mem[830] = 4'b0110;
	mem[831] = 4'b0110;
	mem[832] = 4'b0110;
	mem[833] = 4'b0110;
	mem[834] = 4'b0110;
	mem[835] = 4'b0110;
	mem[836] = 4'b0110;
	mem[837] = 4'b0110;
	mem[838] = 4'b0110;
	mem[839] = 4'b1101;
	mem[840] = 4'b1111;
	mem[841] = 4'b1111;
	mem[842] = 4'b1111;
	mem[843] = 4'b1111;
	mem[844] = 4'b1111;
	mem[845] = 4'b1111;
	mem[846] = 4'b1111;
	mem[847] = 4'b1111;
	mem[848] = 4'b1111;
	mem[849] = 4'b1101;
	mem[850] = 4'b1101;
	mem[851] = 4'b1101;
	mem[852] = 4'b1110;
	mem[853] = 4'b1111;
	mem[854] = 4'b1111;
	mem[855] = 4'b1111;
	mem[856] = 4'b1001;
	mem[857] = 4'b0110;
	mem[858] = 4'b0110;
	mem[859] = 4'b0110;
	mem[860] = 4'b0110;
	mem[861] = 4'b0110;
	mem[862] = 4'b0111;
	mem[863] = 4'b0111;
	mem[864] = 4'b0111;
	mem[865] = 4'b0111;
	mem[866] = 4'b0111;
	mem[867] = 4'b0111;
	mem[868] = 4'b0110;
	mem[869] = 4'b0110;
	mem[870] = 4'b0111;
	mem[871] = 4'b1000;
	mem[872] = 4'b0111;
	mem[873] = 4'b1100;
	mem[874] = 4'b1111;
	mem[875] = 4'b1111;
	mem[876] = 4'b1111;
	mem[877] = 4'b1111;
	mem[878] = 4'b1111;
	mem[879] = 4'b1111;
	mem[880] = 4'b1111;
	mem[881] = 4'b1111;
	mem[882] = 4'b1111;
	mem[883] = 4'b1111;
	mem[884] = 4'b1111;
	mem[885] = 4'b1111;
	mem[886] = 4'b1111;
	mem[887] = 4'b1111;
	mem[888] = 4'b1111;
	mem[889] = 4'b1111;
	mem[890] = 4'b0011;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0111;
	mem[900] = 4'b1100;
	mem[901] = 4'b1101;
	mem[902] = 4'b1101;
	mem[903] = 4'b1101;
	mem[904] = 4'b1101;
	mem[905] = 4'b1101;
	mem[906] = 4'b1101;
	mem[907] = 4'b1101;
	mem[908] = 4'b1101;
	mem[909] = 4'b1101;
	mem[910] = 4'b1101;
	mem[911] = 4'b1101;
	mem[912] = 4'b1101;
	mem[913] = 4'b1101;
	mem[914] = 4'b1101;
	mem[915] = 4'b1101;
	mem[916] = 4'b0111;
	mem[917] = 4'b0101;
	mem[918] = 4'b0101;
	mem[919] = 4'b0101;
	mem[920] = 4'b0101;
	mem[921] = 4'b0101;
	mem[922] = 4'b0101;
	mem[923] = 4'b0110;
	mem[924] = 4'b0110;
	mem[925] = 4'b0110;
	mem[926] = 4'b0110;
	mem[927] = 4'b0110;
	mem[928] = 4'b0101;
	mem[929] = 4'b0101;
	mem[930] = 4'b0101;
	mem[931] = 4'b0110;
	mem[932] = 4'b0110;
	mem[933] = 4'b1101;
	mem[934] = 4'b1111;
	mem[935] = 4'b1111;
	mem[936] = 4'b1111;
	mem[937] = 4'b1111;
	mem[938] = 4'b1111;
	mem[939] = 4'b1111;
	mem[940] = 4'b1111;
	mem[941] = 4'b1111;
	mem[942] = 4'b1111;
	mem[943] = 4'b1111;
	mem[944] = 4'b1111;
	mem[945] = 4'b1111;
	mem[946] = 4'b1111;
	mem[947] = 4'b1111;
	mem[948] = 4'b1111;
	mem[949] = 4'b1111;
	mem[950] = 4'b1010;
	mem[951] = 4'b0110;
	mem[952] = 4'b0110;
	mem[953] = 4'b0110;
	mem[954] = 4'b0110;
	mem[955] = 4'b0110;
	mem[956] = 4'b0110;
	mem[957] = 4'b0110;
	mem[958] = 4'b0110;
	mem[959] = 4'b0110;
	mem[960] = 4'b0110;
	mem[961] = 4'b0110;
	mem[962] = 4'b0110;
	mem[963] = 4'b0110;
	mem[964] = 4'b0110;
	mem[965] = 4'b0110;
	mem[966] = 4'b0110;
	mem[967] = 4'b1101;
	mem[968] = 4'b1111;
	mem[969] = 4'b1111;
	mem[970] = 4'b1111;
	mem[971] = 4'b1111;
	mem[972] = 4'b1111;
	mem[973] = 4'b1111;
	mem[974] = 4'b1111;
	mem[975] = 4'b1111;
	mem[976] = 4'b1110;
	mem[977] = 4'b1101;
	mem[978] = 4'b1101;
	mem[979] = 4'b1110;
	mem[980] = 4'b1111;
	mem[981] = 4'b1111;
	mem[982] = 4'b1111;
	mem[983] = 4'b1111;
	mem[984] = 4'b1000;
	mem[985] = 4'b0110;
	mem[986] = 4'b0110;
	mem[987] = 4'b0110;
	mem[988] = 4'b0110;
	mem[989] = 4'b0110;
	mem[990] = 4'b0110;
	mem[991] = 4'b0111;
	mem[992] = 4'b0111;
	mem[993] = 4'b0111;
	mem[994] = 4'b0111;
	mem[995] = 4'b0111;
	mem[996] = 4'b0111;
	mem[997] = 4'b0111;
	mem[998] = 4'b0111;
	mem[999] = 4'b0101;
	mem[1000] = 4'b0100;
	mem[1001] = 4'b1011;
	mem[1002] = 4'b1111;
	mem[1003] = 4'b1111;
	mem[1004] = 4'b1111;
	mem[1005] = 4'b1111;
	mem[1006] = 4'b1111;
	mem[1007] = 4'b1111;
	mem[1008] = 4'b1111;
	mem[1009] = 4'b1111;
	mem[1010] = 4'b1111;
	mem[1011] = 4'b1111;
	mem[1012] = 4'b1111;
	mem[1013] = 4'b1111;
	mem[1014] = 4'b1111;
	mem[1015] = 4'b1111;
	mem[1016] = 4'b1111;
	mem[1017] = 4'b1111;
	mem[1018] = 4'b0011;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0111;
	mem[1028] = 4'b1100;
	mem[1029] = 4'b1101;
	mem[1030] = 4'b1101;
	mem[1031] = 4'b1101;
	mem[1032] = 4'b1101;
	mem[1033] = 4'b1101;
	mem[1034] = 4'b1101;
	mem[1035] = 4'b1101;
	mem[1036] = 4'b1101;
	mem[1037] = 4'b1101;
	mem[1038] = 4'b1101;
	mem[1039] = 4'b1101;
	mem[1040] = 4'b1101;
	mem[1041] = 4'b1101;
	mem[1042] = 4'b1101;
	mem[1043] = 4'b1101;
	mem[1044] = 4'b0111;
	mem[1045] = 4'b0101;
	mem[1046] = 4'b0101;
	mem[1047] = 4'b0101;
	mem[1048] = 4'b0101;
	mem[1049] = 4'b0101;
	mem[1050] = 4'b0110;
	mem[1051] = 4'b0110;
	mem[1052] = 4'b0110;
	mem[1053] = 4'b0110;
	mem[1054] = 4'b0110;
	mem[1055] = 4'b0101;
	mem[1056] = 4'b0101;
	mem[1057] = 4'b0110;
	mem[1058] = 4'b0111;
	mem[1059] = 4'b0110;
	mem[1060] = 4'b0110;
	mem[1061] = 4'b1100;
	mem[1062] = 4'b1111;
	mem[1063] = 4'b1111;
	mem[1064] = 4'b1111;
	mem[1065] = 4'b1111;
	mem[1066] = 4'b1111;
	mem[1067] = 4'b1111;
	mem[1068] = 4'b1111;
	mem[1069] = 4'b1111;
	mem[1070] = 4'b1111;
	mem[1071] = 4'b1111;
	mem[1072] = 4'b1111;
	mem[1073] = 4'b1111;
	mem[1074] = 4'b1111;
	mem[1075] = 4'b1111;
	mem[1076] = 4'b1111;
	mem[1077] = 4'b1111;
	mem[1078] = 4'b1010;
	mem[1079] = 4'b0110;
	mem[1080] = 4'b0110;
	mem[1081] = 4'b0110;
	mem[1082] = 4'b0110;
	mem[1083] = 4'b0110;
	mem[1084] = 4'b0110;
	mem[1085] = 4'b0110;
	mem[1086] = 4'b0110;
	mem[1087] = 4'b0110;
	mem[1088] = 4'b0110;
	mem[1089] = 4'b0110;
	mem[1090] = 4'b0110;
	mem[1091] = 4'b0110;
	mem[1092] = 4'b0110;
	mem[1093] = 4'b0111;
	mem[1094] = 4'b0111;
	mem[1095] = 4'b1101;
	mem[1096] = 4'b1111;
	mem[1097] = 4'b1111;
	mem[1098] = 4'b1111;
	mem[1099] = 4'b1111;
	mem[1100] = 4'b1111;
	mem[1101] = 4'b1111;
	mem[1102] = 4'b1111;
	mem[1103] = 4'b1111;
	mem[1104] = 4'b1110;
	mem[1105] = 4'b1101;
	mem[1106] = 4'b1101;
	mem[1107] = 4'b1110;
	mem[1108] = 4'b1111;
	mem[1109] = 4'b1111;
	mem[1110] = 4'b1111;
	mem[1111] = 4'b1110;
	mem[1112] = 4'b1000;
	mem[1113] = 4'b0111;
	mem[1114] = 4'b0111;
	mem[1115] = 4'b0110;
	mem[1116] = 4'b0110;
	mem[1117] = 4'b0110;
	mem[1118] = 4'b0110;
	mem[1119] = 4'b0110;
	mem[1120] = 4'b0110;
	mem[1121] = 4'b0101;
	mem[1122] = 4'b0011;
	mem[1123] = 4'b0010;
	mem[1124] = 4'b0001;
	mem[1125] = 4'b0001;
	mem[1126] = 4'b0000;
	mem[1127] = 4'b0000;
	mem[1128] = 4'b0000;
	mem[1129] = 4'b1010;
	mem[1130] = 4'b1111;
	mem[1131] = 4'b1111;
	mem[1132] = 4'b1111;
	mem[1133] = 4'b1111;
	mem[1134] = 4'b1111;
	mem[1135] = 4'b1111;
	mem[1136] = 4'b1111;
	mem[1137] = 4'b1111;
	mem[1138] = 4'b1111;
	mem[1139] = 4'b1111;
	mem[1140] = 4'b1111;
	mem[1141] = 4'b1111;
	mem[1142] = 4'b1111;
	mem[1143] = 4'b1111;
	mem[1144] = 4'b1111;
	mem[1145] = 4'b1111;
	mem[1146] = 4'b0011;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0111;
	mem[1156] = 4'b1100;
	mem[1157] = 4'b1101;
	mem[1158] = 4'b1101;
	mem[1159] = 4'b1101;
	mem[1160] = 4'b1101;
	mem[1161] = 4'b1101;
	mem[1162] = 4'b1101;
	mem[1163] = 4'b1101;
	mem[1164] = 4'b1101;
	mem[1165] = 4'b1101;
	mem[1166] = 4'b1101;
	mem[1167] = 4'b1101;
	mem[1168] = 4'b1101;
	mem[1169] = 4'b1101;
	mem[1170] = 4'b1101;
	mem[1171] = 4'b1101;
	mem[1172] = 4'b0111;
	mem[1173] = 4'b0101;
	mem[1174] = 4'b0101;
	mem[1175] = 4'b0101;
	mem[1176] = 4'b0110;
	mem[1177] = 4'b0110;
	mem[1178] = 4'b0110;
	mem[1179] = 4'b0110;
	mem[1180] = 4'b0110;
	mem[1181] = 4'b0110;
	mem[1182] = 4'b0101;
	mem[1183] = 4'b0101;
	mem[1184] = 4'b0110;
	mem[1185] = 4'b0110;
	mem[1186] = 4'b0110;
	mem[1187] = 4'b0101;
	mem[1188] = 4'b0101;
	mem[1189] = 4'b1011;
	mem[1190] = 4'b1101;
	mem[1191] = 4'b1111;
	mem[1192] = 4'b1111;
	mem[1193] = 4'b1111;
	mem[1194] = 4'b1111;
	mem[1195] = 4'b1111;
	mem[1196] = 4'b1111;
	mem[1197] = 4'b1111;
	mem[1198] = 4'b1111;
	mem[1199] = 4'b1111;
	mem[1200] = 4'b1111;
	mem[1201] = 4'b1111;
	mem[1202] = 4'b1111;
	mem[1203] = 4'b1111;
	mem[1204] = 4'b1111;
	mem[1205] = 4'b1111;
	mem[1206] = 4'b1010;
	mem[1207] = 4'b0110;
	mem[1208] = 4'b0110;
	mem[1209] = 4'b0110;
	mem[1210] = 4'b0110;
	mem[1211] = 4'b0110;
	mem[1212] = 4'b0110;
	mem[1213] = 4'b0110;
	mem[1214] = 4'b0110;
	mem[1215] = 4'b0110;
	mem[1216] = 4'b0110;
	mem[1217] = 4'b0110;
	mem[1218] = 4'b0110;
	mem[1219] = 4'b0111;
	mem[1220] = 4'b0111;
	mem[1221] = 4'b0111;
	mem[1222] = 4'b0111;
	mem[1223] = 4'b1101;
	mem[1224] = 4'b1111;
	mem[1225] = 4'b1111;
	mem[1226] = 4'b1111;
	mem[1227] = 4'b1111;
	mem[1228] = 4'b1111;
	mem[1229] = 4'b1111;
	mem[1230] = 4'b1111;
	mem[1231] = 4'b1111;
	mem[1232] = 4'b1110;
	mem[1233] = 4'b1101;
	mem[1234] = 4'b1101;
	mem[1235] = 4'b1110;
	mem[1236] = 4'b1111;
	mem[1237] = 4'b1111;
	mem[1238] = 4'b1110;
	mem[1239] = 4'b1101;
	mem[1240] = 4'b1000;
	mem[1241] = 4'b1000;
	mem[1242] = 4'b0111;
	mem[1243] = 4'b0101;
	mem[1244] = 4'b0011;
	mem[1245] = 4'b0010;
	mem[1246] = 4'b0001;
	mem[1247] = 4'b0000;
	mem[1248] = 4'b0000;
	mem[1249] = 4'b0000;
	mem[1250] = 4'b0000;
	mem[1251] = 4'b0000;
	mem[1252] = 4'b0000;
	mem[1253] = 4'b0000;
	mem[1254] = 4'b0000;
	mem[1255] = 4'b0000;
	mem[1256] = 4'b0000;
	mem[1257] = 4'b1010;
	mem[1258] = 4'b1111;
	mem[1259] = 4'b1111;
	mem[1260] = 4'b1111;
	mem[1261] = 4'b1111;
	mem[1262] = 4'b1111;
	mem[1263] = 4'b1111;
	mem[1264] = 4'b1111;
	mem[1265] = 4'b1111;
	mem[1266] = 4'b1111;
	mem[1267] = 4'b1111;
	mem[1268] = 4'b1111;
	mem[1269] = 4'b1111;
	mem[1270] = 4'b1111;
	mem[1271] = 4'b1111;
	mem[1272] = 4'b1111;
	mem[1273] = 4'b1111;
	mem[1274] = 4'b0011;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0111;
	mem[1284] = 4'b1100;
	mem[1285] = 4'b1101;
	mem[1286] = 4'b1101;
	mem[1287] = 4'b1101;
	mem[1288] = 4'b1101;
	mem[1289] = 4'b1101;
	mem[1290] = 4'b1101;
	mem[1291] = 4'b1101;
	mem[1292] = 4'b1101;
	mem[1293] = 4'b1101;
	mem[1294] = 4'b1101;
	mem[1295] = 4'b1101;
	mem[1296] = 4'b1101;
	mem[1297] = 4'b1101;
	mem[1298] = 4'b1101;
	mem[1299] = 4'b1101;
	mem[1300] = 4'b0111;
	mem[1301] = 4'b0101;
	mem[1302] = 4'b0110;
	mem[1303] = 4'b0110;
	mem[1304] = 4'b0110;
	mem[1305] = 4'b0110;
	mem[1306] = 4'b0110;
	mem[1307] = 4'b0110;
	mem[1308] = 4'b0110;
	mem[1309] = 4'b0110;
	mem[1310] = 4'b0110;
	mem[1311] = 4'b0101;
	mem[1312] = 4'b0110;
	mem[1313] = 4'b0110;
	mem[1314] = 4'b0101;
	mem[1315] = 4'b0101;
	mem[1316] = 4'b0110;
	mem[1317] = 4'b1100;
	mem[1318] = 4'b1101;
	mem[1319] = 4'b1110;
	mem[1320] = 4'b1111;
	mem[1321] = 4'b1111;
	mem[1322] = 4'b1111;
	mem[1323] = 4'b1111;
	mem[1324] = 4'b1111;
	mem[1325] = 4'b1111;
	mem[1326] = 4'b1111;
	mem[1327] = 4'b1111;
	mem[1328] = 4'b1111;
	mem[1329] = 4'b1111;
	mem[1330] = 4'b1111;
	mem[1331] = 4'b1111;
	mem[1332] = 4'b1111;
	mem[1333] = 4'b1111;
	mem[1334] = 4'b1010;
	mem[1335] = 4'b0110;
	mem[1336] = 4'b0110;
	mem[1337] = 4'b0110;
	mem[1338] = 4'b0110;
	mem[1339] = 4'b0110;
	mem[1340] = 4'b0110;
	mem[1341] = 4'b0110;
	mem[1342] = 4'b0110;
	mem[1343] = 4'b0110;
	mem[1344] = 4'b0110;
	mem[1345] = 4'b0111;
	mem[1346] = 4'b0111;
	mem[1347] = 4'b0111;
	mem[1348] = 4'b0111;
	mem[1349] = 4'b0111;
	mem[1350] = 4'b0111;
	mem[1351] = 4'b1101;
	mem[1352] = 4'b1111;
	mem[1353] = 4'b1111;
	mem[1354] = 4'b1111;
	mem[1355] = 4'b1111;
	mem[1356] = 4'b1111;
	mem[1357] = 4'b1111;
	mem[1358] = 4'b1111;
	mem[1359] = 4'b1111;
	mem[1360] = 4'b1111;
	mem[1361] = 4'b1101;
	mem[1362] = 4'b1110;
	mem[1363] = 4'b1111;
	mem[1364] = 4'b1111;
	mem[1365] = 4'b1111;
	mem[1366] = 4'b1101;
	mem[1367] = 4'b1101;
	mem[1368] = 4'b0101;
	mem[1369] = 4'b0001;
	mem[1370] = 4'b0000;
	mem[1371] = 4'b0000;
	mem[1372] = 4'b0000;
	mem[1373] = 4'b0000;
	mem[1374] = 4'b0000;
	mem[1375] = 4'b0000;
	mem[1376] = 4'b0000;
	mem[1377] = 4'b0000;
	mem[1378] = 4'b0001;
	mem[1379] = 4'b0000;
	mem[1380] = 4'b0000;
	mem[1381] = 4'b0000;
	mem[1382] = 4'b0000;
	mem[1383] = 4'b0000;
	mem[1384] = 4'b0000;
	mem[1385] = 4'b1010;
	mem[1386] = 4'b1111;
	mem[1387] = 4'b1111;
	mem[1388] = 4'b1111;
	mem[1389] = 4'b1111;
	mem[1390] = 4'b1111;
	mem[1391] = 4'b1111;
	mem[1392] = 4'b1111;
	mem[1393] = 4'b1111;
	mem[1394] = 4'b1111;
	mem[1395] = 4'b1111;
	mem[1396] = 4'b1111;
	mem[1397] = 4'b1111;
	mem[1398] = 4'b1111;
	mem[1399] = 4'b1111;
	mem[1400] = 4'b1111;
	mem[1401] = 4'b1111;
	mem[1402] = 4'b0011;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0111;
	mem[1412] = 4'b1100;
	mem[1413] = 4'b1101;
	mem[1414] = 4'b1101;
	mem[1415] = 4'b1101;
	mem[1416] = 4'b1101;
	mem[1417] = 4'b1101;
	mem[1418] = 4'b1101;
	mem[1419] = 4'b1101;
	mem[1420] = 4'b1101;
	mem[1421] = 4'b1101;
	mem[1422] = 4'b1101;
	mem[1423] = 4'b1101;
	mem[1424] = 4'b1101;
	mem[1425] = 4'b1101;
	mem[1426] = 4'b1101;
	mem[1427] = 4'b1101;
	mem[1428] = 4'b1000;
	mem[1429] = 4'b0110;
	mem[1430] = 4'b0110;
	mem[1431] = 4'b0110;
	mem[1432] = 4'b0110;
	mem[1433] = 4'b0110;
	mem[1434] = 4'b0110;
	mem[1435] = 4'b0110;
	mem[1436] = 4'b0110;
	mem[1437] = 4'b0110;
	mem[1438] = 4'b0110;
	mem[1439] = 4'b0101;
	mem[1440] = 4'b0101;
	mem[1441] = 4'b0101;
	mem[1442] = 4'b0101;
	mem[1443] = 4'b0110;
	mem[1444] = 4'b0111;
	mem[1445] = 4'b1101;
	mem[1446] = 4'b1101;
	mem[1447] = 4'b1110;
	mem[1448] = 4'b1111;
	mem[1449] = 4'b1111;
	mem[1450] = 4'b1111;
	mem[1451] = 4'b1111;
	mem[1452] = 4'b1111;
	mem[1453] = 4'b1111;
	mem[1454] = 4'b1111;
	mem[1455] = 4'b1111;
	mem[1456] = 4'b1111;
	mem[1457] = 4'b1111;
	mem[1458] = 4'b1111;
	mem[1459] = 4'b1111;
	mem[1460] = 4'b1111;
	mem[1461] = 4'b1111;
	mem[1462] = 4'b1010;
	mem[1463] = 4'b0110;
	mem[1464] = 4'b0110;
	mem[1465] = 4'b0110;
	mem[1466] = 4'b0110;
	mem[1467] = 4'b0110;
	mem[1468] = 4'b0110;
	mem[1469] = 4'b0110;
	mem[1470] = 4'b0110;
	mem[1471] = 4'b0111;
	mem[1472] = 4'b0111;
	mem[1473] = 4'b0111;
	mem[1474] = 4'b0111;
	mem[1475] = 4'b0111;
	mem[1476] = 4'b0111;
	mem[1477] = 4'b0111;
	mem[1478] = 4'b0111;
	mem[1479] = 4'b1101;
	mem[1480] = 4'b1111;
	mem[1481] = 4'b1111;
	mem[1482] = 4'b1111;
	mem[1483] = 4'b1111;
	mem[1484] = 4'b1111;
	mem[1485] = 4'b1111;
	mem[1486] = 4'b1111;
	mem[1487] = 4'b1111;
	mem[1488] = 4'b1111;
	mem[1489] = 4'b1111;
	mem[1490] = 4'b1111;
	mem[1491] = 4'b1111;
	mem[1492] = 4'b1111;
	mem[1493] = 4'b1110;
	mem[1494] = 4'b1101;
	mem[1495] = 4'b1101;
	mem[1496] = 4'b0101;
	mem[1497] = 4'b0000;
	mem[1498] = 4'b0000;
	mem[1499] = 4'b0000;
	mem[1500] = 4'b0000;
	mem[1501] = 4'b0000;
	mem[1502] = 4'b0000;
	mem[1503] = 4'b0000;
	mem[1504] = 4'b0000;
	mem[1505] = 4'b0001;
	mem[1506] = 4'b0000;
	mem[1507] = 4'b0000;
	mem[1508] = 4'b0000;
	mem[1509] = 4'b0000;
	mem[1510] = 4'b0000;
	mem[1511] = 4'b0000;
	mem[1512] = 4'b0000;
	mem[1513] = 4'b1010;
	mem[1514] = 4'b1111;
	mem[1515] = 4'b1111;
	mem[1516] = 4'b1111;
	mem[1517] = 4'b1111;
	mem[1518] = 4'b1111;
	mem[1519] = 4'b1111;
	mem[1520] = 4'b1111;
	mem[1521] = 4'b1111;
	mem[1522] = 4'b1111;
	mem[1523] = 4'b1111;
	mem[1524] = 4'b1111;
	mem[1525] = 4'b1111;
	mem[1526] = 4'b1111;
	mem[1527] = 4'b1111;
	mem[1528] = 4'b1111;
	mem[1529] = 4'b1111;
	mem[1530] = 4'b0011;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0111;
	mem[1540] = 4'b1100;
	mem[1541] = 4'b1101;
	mem[1542] = 4'b1101;
	mem[1543] = 4'b1101;
	mem[1544] = 4'b1101;
	mem[1545] = 4'b1101;
	mem[1546] = 4'b1101;
	mem[1547] = 4'b1101;
	mem[1548] = 4'b1101;
	mem[1549] = 4'b1101;
	mem[1550] = 4'b1101;
	mem[1551] = 4'b1101;
	mem[1552] = 4'b1101;
	mem[1553] = 4'b1101;
	mem[1554] = 4'b1101;
	mem[1555] = 4'b1101;
	mem[1556] = 4'b1000;
	mem[1557] = 4'b0110;
	mem[1558] = 4'b0110;
	mem[1559] = 4'b0110;
	mem[1560] = 4'b0110;
	mem[1561] = 4'b0110;
	mem[1562] = 4'b0110;
	mem[1563] = 4'b0110;
	mem[1564] = 4'b0110;
	mem[1565] = 4'b0110;
	mem[1566] = 4'b0110;
	mem[1567] = 4'b0110;
	mem[1568] = 4'b0110;
	mem[1569] = 4'b0110;
	mem[1570] = 4'b0111;
	mem[1571] = 4'b0111;
	mem[1572] = 4'b0110;
	mem[1573] = 4'b1100;
	mem[1574] = 4'b1101;
	mem[1575] = 4'b1111;
	mem[1576] = 4'b1111;
	mem[1577] = 4'b1111;
	mem[1578] = 4'b1111;
	mem[1579] = 4'b1111;
	mem[1580] = 4'b1111;
	mem[1581] = 4'b1111;
	mem[1582] = 4'b1111;
	mem[1583] = 4'b1111;
	mem[1584] = 4'b1111;
	mem[1585] = 4'b1111;
	mem[1586] = 4'b1111;
	mem[1587] = 4'b1111;
	mem[1588] = 4'b1111;
	mem[1589] = 4'b1111;
	mem[1590] = 4'b1010;
	mem[1591] = 4'b0110;
	mem[1592] = 4'b0110;
	mem[1593] = 4'b0110;
	mem[1594] = 4'b0110;
	mem[1595] = 4'b0110;
	mem[1596] = 4'b0110;
	mem[1597] = 4'b0111;
	mem[1598] = 4'b0111;
	mem[1599] = 4'b0111;
	mem[1600] = 4'b0111;
	mem[1601] = 4'b0111;
	mem[1602] = 4'b0111;
	mem[1603] = 4'b0111;
	mem[1604] = 4'b0111;
	mem[1605] = 4'b0111;
	mem[1606] = 4'b0111;
	mem[1607] = 4'b1101;
	mem[1608] = 4'b1111;
	mem[1609] = 4'b1111;
	mem[1610] = 4'b1111;
	mem[1611] = 4'b1111;
	mem[1612] = 4'b1111;
	mem[1613] = 4'b1111;
	mem[1614] = 4'b1111;
	mem[1615] = 4'b1111;
	mem[1616] = 4'b1111;
	mem[1617] = 4'b1111;
	mem[1618] = 4'b1111;
	mem[1619] = 4'b1111;
	mem[1620] = 4'b1111;
	mem[1621] = 4'b1101;
	mem[1622] = 4'b1101;
	mem[1623] = 4'b1110;
	mem[1624] = 4'b0100;
	mem[1625] = 4'b0000;
	mem[1626] = 4'b0000;
	mem[1627] = 4'b0000;
	mem[1628] = 4'b0000;
	mem[1629] = 4'b0000;
	mem[1630] = 4'b0001;
	mem[1631] = 4'b0001;
	mem[1632] = 4'b0001;
	mem[1633] = 4'b0000;
	mem[1634] = 4'b0000;
	mem[1635] = 4'b0000;
	mem[1636] = 4'b0000;
	mem[1637] = 4'b0000;
	mem[1638] = 4'b0000;
	mem[1639] = 4'b0000;
	mem[1640] = 4'b0000;
	mem[1641] = 4'b1010;
	mem[1642] = 4'b1111;
	mem[1643] = 4'b1111;
	mem[1644] = 4'b1111;
	mem[1645] = 4'b1111;
	mem[1646] = 4'b1111;
	mem[1647] = 4'b1111;
	mem[1648] = 4'b1111;
	mem[1649] = 4'b1111;
	mem[1650] = 4'b1111;
	mem[1651] = 4'b1111;
	mem[1652] = 4'b1111;
	mem[1653] = 4'b1111;
	mem[1654] = 4'b1111;
	mem[1655] = 4'b1111;
	mem[1656] = 4'b1111;
	mem[1657] = 4'b1111;
	mem[1658] = 4'b0011;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0111;
	mem[1668] = 4'b1100;
	mem[1669] = 4'b1101;
	mem[1670] = 4'b1101;
	mem[1671] = 4'b1101;
	mem[1672] = 4'b1101;
	mem[1673] = 4'b1101;
	mem[1674] = 4'b1101;
	mem[1675] = 4'b1101;
	mem[1676] = 4'b1101;
	mem[1677] = 4'b1101;
	mem[1678] = 4'b1101;
	mem[1679] = 4'b1101;
	mem[1680] = 4'b1101;
	mem[1681] = 4'b1101;
	mem[1682] = 4'b1101;
	mem[1683] = 4'b1101;
	mem[1684] = 4'b1000;
	mem[1685] = 4'b0110;
	mem[1686] = 4'b0110;
	mem[1687] = 4'b0110;
	mem[1688] = 4'b0110;
	mem[1689] = 4'b0110;
	mem[1690] = 4'b0101;
	mem[1691] = 4'b0101;
	mem[1692] = 4'b0101;
	mem[1693] = 4'b0110;
	mem[1694] = 4'b0110;
	mem[1695] = 4'b0110;
	mem[1696] = 4'b0110;
	mem[1697] = 4'b0110;
	mem[1698] = 4'b0110;
	mem[1699] = 4'b0110;
	mem[1700] = 4'b0110;
	mem[1701] = 4'b1011;
	mem[1702] = 4'b1110;
	mem[1703] = 4'b1111;
	mem[1704] = 4'b1111;
	mem[1705] = 4'b1111;
	mem[1706] = 4'b1111;
	mem[1707] = 4'b1111;
	mem[1708] = 4'b1111;
	mem[1709] = 4'b1111;
	mem[1710] = 4'b1111;
	mem[1711] = 4'b1111;
	mem[1712] = 4'b1111;
	mem[1713] = 4'b1111;
	mem[1714] = 4'b1111;
	mem[1715] = 4'b1111;
	mem[1716] = 4'b1111;
	mem[1717] = 4'b1111;
	mem[1718] = 4'b1010;
	mem[1719] = 4'b0110;
	mem[1720] = 4'b0110;
	mem[1721] = 4'b0110;
	mem[1722] = 4'b0110;
	mem[1723] = 4'b0110;
	mem[1724] = 4'b0111;
	mem[1725] = 4'b0111;
	mem[1726] = 4'b0111;
	mem[1727] = 4'b0111;
	mem[1728] = 4'b0111;
	mem[1729] = 4'b0111;
	mem[1730] = 4'b0111;
	mem[1731] = 4'b0111;
	mem[1732] = 4'b0111;
	mem[1733] = 4'b0111;
	mem[1734] = 4'b0111;
	mem[1735] = 4'b1101;
	mem[1736] = 4'b1111;
	mem[1737] = 4'b1111;
	mem[1738] = 4'b1111;
	mem[1739] = 4'b1111;
	mem[1740] = 4'b1111;
	mem[1741] = 4'b1111;
	mem[1742] = 4'b1111;
	mem[1743] = 4'b1111;
	mem[1744] = 4'b1111;
	mem[1745] = 4'b1111;
	mem[1746] = 4'b1111;
	mem[1747] = 4'b1111;
	mem[1748] = 4'b1110;
	mem[1749] = 4'b1101;
	mem[1750] = 4'b1101;
	mem[1751] = 4'b1101;
	mem[1752] = 4'b0100;
	mem[1753] = 4'b0000;
	mem[1754] = 4'b0000;
	mem[1755] = 4'b0000;
	mem[1756] = 4'b0000;
	mem[1757] = 4'b0000;
	mem[1758] = 4'b0001;
	mem[1759] = 4'b0000;
	mem[1760] = 4'b0000;
	mem[1761] = 4'b0000;
	mem[1762] = 4'b0000;
	mem[1763] = 4'b0000;
	mem[1764] = 4'b0000;
	mem[1765] = 4'b0000;
	mem[1766] = 4'b0000;
	mem[1767] = 4'b0000;
	mem[1768] = 4'b0000;
	mem[1769] = 4'b1010;
	mem[1770] = 4'b1111;
	mem[1771] = 4'b1111;
	mem[1772] = 4'b1111;
	mem[1773] = 4'b1111;
	mem[1774] = 4'b1111;
	mem[1775] = 4'b1111;
	mem[1776] = 4'b1111;
	mem[1777] = 4'b1111;
	mem[1778] = 4'b1111;
	mem[1779] = 4'b1111;
	mem[1780] = 4'b1111;
	mem[1781] = 4'b1111;
	mem[1782] = 4'b1111;
	mem[1783] = 4'b1111;
	mem[1784] = 4'b1111;
	mem[1785] = 4'b1111;
	mem[1786] = 4'b0011;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0111;
	mem[1796] = 4'b1100;
	mem[1797] = 4'b1101;
	mem[1798] = 4'b1101;
	mem[1799] = 4'b1101;
	mem[1800] = 4'b1101;
	mem[1801] = 4'b1101;
	mem[1802] = 4'b1101;
	mem[1803] = 4'b1101;
	mem[1804] = 4'b1101;
	mem[1805] = 4'b1101;
	mem[1806] = 4'b1101;
	mem[1807] = 4'b1101;
	mem[1808] = 4'b1101;
	mem[1809] = 4'b1101;
	mem[1810] = 4'b1101;
	mem[1811] = 4'b1101;
	mem[1812] = 4'b1000;
	mem[1813] = 4'b0110;
	mem[1814] = 4'b0110;
	mem[1815] = 4'b0110;
	mem[1816] = 4'b0110;
	mem[1817] = 4'b0101;
	mem[1818] = 4'b0101;
	mem[1819] = 4'b0101;
	mem[1820] = 4'b0101;
	mem[1821] = 4'b0101;
	mem[1822] = 4'b0110;
	mem[1823] = 4'b0110;
	mem[1824] = 4'b0110;
	mem[1825] = 4'b0110;
	mem[1826] = 4'b0101;
	mem[1827] = 4'b0101;
	mem[1828] = 4'b0101;
	mem[1829] = 4'b1100;
	mem[1830] = 4'b1111;
	mem[1831] = 4'b1111;
	mem[1832] = 4'b1111;
	mem[1833] = 4'b1111;
	mem[1834] = 4'b1111;
	mem[1835] = 4'b1111;
	mem[1836] = 4'b1111;
	mem[1837] = 4'b1111;
	mem[1838] = 4'b1111;
	mem[1839] = 4'b1111;
	mem[1840] = 4'b1111;
	mem[1841] = 4'b1111;
	mem[1842] = 4'b1111;
	mem[1843] = 4'b1111;
	mem[1844] = 4'b1111;
	mem[1845] = 4'b1111;
	mem[1846] = 4'b1010;
	mem[1847] = 4'b0110;
	mem[1848] = 4'b0110;
	mem[1849] = 4'b0110;
	mem[1850] = 4'b0111;
	mem[1851] = 4'b0111;
	mem[1852] = 4'b0111;
	mem[1853] = 4'b0111;
	mem[1854] = 4'b0111;
	mem[1855] = 4'b0111;
	mem[1856] = 4'b0111;
	mem[1857] = 4'b0111;
	mem[1858] = 4'b0111;
	mem[1859] = 4'b0111;
	mem[1860] = 4'b0111;
	mem[1861] = 4'b0101;
	mem[1862] = 4'b0011;
	mem[1863] = 4'b1100;
	mem[1864] = 4'b1111;
	mem[1865] = 4'b1111;
	mem[1866] = 4'b1111;
	mem[1867] = 4'b1111;
	mem[1868] = 4'b1111;
	mem[1869] = 4'b1111;
	mem[1870] = 4'b1111;
	mem[1871] = 4'b1111;
	mem[1872] = 4'b1111;
	mem[1873] = 4'b1111;
	mem[1874] = 4'b1111;
	mem[1875] = 4'b1111;
	mem[1876] = 4'b1111;
	mem[1877] = 4'b1101;
	mem[1878] = 4'b1101;
	mem[1879] = 4'b1101;
	mem[1880] = 4'b0100;
	mem[1881] = 4'b0000;
	mem[1882] = 4'b0000;
	mem[1883] = 4'b0000;
	mem[1884] = 4'b0000;
	mem[1885] = 4'b0000;
	mem[1886] = 4'b0001;
	mem[1887] = 4'b0000;
	mem[1888] = 4'b0000;
	mem[1889] = 4'b0000;
	mem[1890] = 4'b0000;
	mem[1891] = 4'b0000;
	mem[1892] = 4'b0000;
	mem[1893] = 4'b0000;
	mem[1894] = 4'b0000;
	mem[1895] = 4'b0000;
	mem[1896] = 4'b0000;
	mem[1897] = 4'b1010;
	mem[1898] = 4'b1111;
	mem[1899] = 4'b1111;
	mem[1900] = 4'b1111;
	mem[1901] = 4'b1111;
	mem[1902] = 4'b1111;
	mem[1903] = 4'b1111;
	mem[1904] = 4'b1111;
	mem[1905] = 4'b1111;
	mem[1906] = 4'b1111;
	mem[1907] = 4'b1111;
	mem[1908] = 4'b1111;
	mem[1909] = 4'b1111;
	mem[1910] = 4'b1111;
	mem[1911] = 4'b1111;
	mem[1912] = 4'b1111;
	mem[1913] = 4'b1111;
	mem[1914] = 4'b0011;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0111;
	mem[1924] = 4'b1100;
	mem[1925] = 4'b1101;
	mem[1926] = 4'b1101;
	mem[1927] = 4'b1101;
	mem[1928] = 4'b1101;
	mem[1929] = 4'b1101;
	mem[1930] = 4'b1101;
	mem[1931] = 4'b1101;
	mem[1932] = 4'b1101;
	mem[1933] = 4'b1101;
	mem[1934] = 4'b1101;
	mem[1935] = 4'b1101;
	mem[1936] = 4'b1101;
	mem[1937] = 4'b1101;
	mem[1938] = 4'b1101;
	mem[1939] = 4'b1110;
	mem[1940] = 4'b1000;
	mem[1941] = 4'b0110;
	mem[1942] = 4'b0110;
	mem[1943] = 4'b0110;
	mem[1944] = 4'b0110;
	mem[1945] = 4'b0101;
	mem[1946] = 4'b0110;
	mem[1947] = 4'b0111;
	mem[1948] = 4'b0110;
	mem[1949] = 4'b0101;
	mem[1950] = 4'b0101;
	mem[1951] = 4'b0110;
	mem[1952] = 4'b0110;
	mem[1953] = 4'b0110;
	mem[1954] = 4'b0110;
	mem[1955] = 4'b0111;
	mem[1956] = 4'b0111;
	mem[1957] = 4'b1101;
	mem[1958] = 4'b1111;
	mem[1959] = 4'b1111;
	mem[1960] = 4'b1111;
	mem[1961] = 4'b1111;
	mem[1962] = 4'b1111;
	mem[1963] = 4'b1111;
	mem[1964] = 4'b1111;
	mem[1965] = 4'b1111;
	mem[1966] = 4'b1111;
	mem[1967] = 4'b1111;
	mem[1968] = 4'b1111;
	mem[1969] = 4'b1111;
	mem[1970] = 4'b1111;
	mem[1971] = 4'b1111;
	mem[1972] = 4'b1111;
	mem[1973] = 4'b1111;
	mem[1974] = 4'b1010;
	mem[1975] = 4'b0110;
	mem[1976] = 4'b0111;
	mem[1977] = 4'b0111;
	mem[1978] = 4'b0111;
	mem[1979] = 4'b0111;
	mem[1980] = 4'b0111;
	mem[1981] = 4'b0111;
	mem[1982] = 4'b0111;
	mem[1983] = 4'b0111;
	mem[1984] = 4'b0110;
	mem[1985] = 4'b0110;
	mem[1986] = 4'b0100;
	mem[1987] = 4'b0010;
	mem[1988] = 4'b0000;
	mem[1989] = 4'b0000;
	mem[1990] = 4'b0000;
	mem[1991] = 4'b1100;
	mem[1992] = 4'b1111;
	mem[1993] = 4'b1111;
	mem[1994] = 4'b1111;
	mem[1995] = 4'b1111;
	mem[1996] = 4'b1111;
	mem[1997] = 4'b1111;
	mem[1998] = 4'b1111;
	mem[1999] = 4'b1111;
	mem[2000] = 4'b1111;
	mem[2001] = 4'b1111;
	mem[2002] = 4'b1111;
	mem[2003] = 4'b1111;
	mem[2004] = 4'b1111;
	mem[2005] = 4'b1101;
	mem[2006] = 4'b1101;
	mem[2007] = 4'b1101;
	mem[2008] = 4'b0011;
	mem[2009] = 4'b0000;
	mem[2010] = 4'b0000;
	mem[2011] = 4'b0000;
	mem[2012] = 4'b0000;
	mem[2013] = 4'b0001;
	mem[2014] = 4'b0000;
	mem[2015] = 4'b0000;
	mem[2016] = 4'b0000;
	mem[2017] = 4'b0000;
	mem[2018] = 4'b0000;
	mem[2019] = 4'b0000;
	mem[2020] = 4'b0000;
	mem[2021] = 4'b0000;
	mem[2022] = 4'b0000;
	mem[2023] = 4'b0000;
	mem[2024] = 4'b0000;
	mem[2025] = 4'b1010;
	mem[2026] = 4'b1111;
	mem[2027] = 4'b1111;
	mem[2028] = 4'b1111;
	mem[2029] = 4'b1111;
	mem[2030] = 4'b1111;
	mem[2031] = 4'b1111;
	mem[2032] = 4'b1111;
	mem[2033] = 4'b1111;
	mem[2034] = 4'b1111;
	mem[2035] = 4'b1111;
	mem[2036] = 4'b1111;
	mem[2037] = 4'b1111;
	mem[2038] = 4'b1111;
	mem[2039] = 4'b1111;
	mem[2040] = 4'b1111;
	mem[2041] = 4'b1111;
	mem[2042] = 4'b0011;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0111;
	mem[2052] = 4'b1100;
	mem[2053] = 4'b1101;
	mem[2054] = 4'b1101;
	mem[2055] = 4'b1101;
	mem[2056] = 4'b1101;
	mem[2057] = 4'b1101;
	mem[2058] = 4'b1101;
	mem[2059] = 4'b1101;
	mem[2060] = 4'b1101;
	mem[2061] = 4'b1101;
	mem[2062] = 4'b1101;
	mem[2063] = 4'b1101;
	mem[2064] = 4'b1101;
	mem[2065] = 4'b1101;
	mem[2066] = 4'b1110;
	mem[2067] = 4'b1110;
	mem[2068] = 4'b1000;
	mem[2069] = 4'b0110;
	mem[2070] = 4'b0110;
	mem[2071] = 4'b0110;
	mem[2072] = 4'b0110;
	mem[2073] = 4'b0101;
	mem[2074] = 4'b0111;
	mem[2075] = 4'b0110;
	mem[2076] = 4'b0110;
	mem[2077] = 4'b0110;
	mem[2078] = 4'b0101;
	mem[2079] = 4'b0101;
	mem[2080] = 4'b0110;
	mem[2081] = 4'b0110;
	mem[2082] = 4'b0110;
	mem[2083] = 4'b0110;
	mem[2084] = 4'b0110;
	mem[2085] = 4'b1101;
	mem[2086] = 4'b1111;
	mem[2087] = 4'b1111;
	mem[2088] = 4'b1111;
	mem[2089] = 4'b1111;
	mem[2090] = 4'b1111;
	mem[2091] = 4'b1111;
	mem[2092] = 4'b1111;
	mem[2093] = 4'b1111;
	mem[2094] = 4'b1111;
	mem[2095] = 4'b1111;
	mem[2096] = 4'b1111;
	mem[2097] = 4'b1111;
	mem[2098] = 4'b1111;
	mem[2099] = 4'b1111;
	mem[2100] = 4'b1111;
	mem[2101] = 4'b1111;
	mem[2102] = 4'b1010;
	mem[2103] = 4'b0111;
	mem[2104] = 4'b0111;
	mem[2105] = 4'b0111;
	mem[2106] = 4'b0111;
	mem[2107] = 4'b0111;
	mem[2108] = 4'b0111;
	mem[2109] = 4'b0111;
	mem[2110] = 4'b0110;
	mem[2111] = 4'b0011;
	mem[2112] = 4'b0001;
	mem[2113] = 4'b0000;
	mem[2114] = 4'b0000;
	mem[2115] = 4'b0000;
	mem[2116] = 4'b0000;
	mem[2117] = 4'b0000;
	mem[2118] = 4'b0000;
	mem[2119] = 4'b1100;
	mem[2120] = 4'b1111;
	mem[2121] = 4'b1111;
	mem[2122] = 4'b1111;
	mem[2123] = 4'b1111;
	mem[2124] = 4'b1111;
	mem[2125] = 4'b1111;
	mem[2126] = 4'b1111;
	mem[2127] = 4'b1111;
	mem[2128] = 4'b1111;
	mem[2129] = 4'b1111;
	mem[2130] = 4'b1111;
	mem[2131] = 4'b1111;
	mem[2132] = 4'b1111;
	mem[2133] = 4'b1111;
	mem[2134] = 4'b1101;
	mem[2135] = 4'b1101;
	mem[2136] = 4'b0011;
	mem[2137] = 4'b0000;
	mem[2138] = 4'b0000;
	mem[2139] = 4'b0000;
	mem[2140] = 4'b0001;
	mem[2141] = 4'b0001;
	mem[2142] = 4'b0000;
	mem[2143] = 4'b0000;
	mem[2144] = 4'b0000;
	mem[2145] = 4'b0000;
	mem[2146] = 4'b0000;
	mem[2147] = 4'b0000;
	mem[2148] = 4'b0000;
	mem[2149] = 4'b0000;
	mem[2150] = 4'b0000;
	mem[2151] = 4'b0000;
	mem[2152] = 4'b0000;
	mem[2153] = 4'b1010;
	mem[2154] = 4'b1111;
	mem[2155] = 4'b1111;
	mem[2156] = 4'b1111;
	mem[2157] = 4'b1111;
	mem[2158] = 4'b1111;
	mem[2159] = 4'b1111;
	mem[2160] = 4'b1111;
	mem[2161] = 4'b1111;
	mem[2162] = 4'b1111;
	mem[2163] = 4'b1111;
	mem[2164] = 4'b1111;
	mem[2165] = 4'b1111;
	mem[2166] = 4'b1111;
	mem[2167] = 4'b1111;
	mem[2168] = 4'b1111;
	mem[2169] = 4'b1111;
	mem[2170] = 4'b0011;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0111;
	mem[2180] = 4'b1100;
	mem[2181] = 4'b1101;
	mem[2182] = 4'b1101;
	mem[2183] = 4'b1101;
	mem[2184] = 4'b1101;
	mem[2185] = 4'b1101;
	mem[2186] = 4'b1101;
	mem[2187] = 4'b1101;
	mem[2188] = 4'b1101;
	mem[2189] = 4'b1101;
	mem[2190] = 4'b1101;
	mem[2191] = 4'b1101;
	mem[2192] = 4'b1110;
	mem[2193] = 4'b1110;
	mem[2194] = 4'b1110;
	mem[2195] = 4'b1110;
	mem[2196] = 4'b1000;
	mem[2197] = 4'b0110;
	mem[2198] = 4'b0110;
	mem[2199] = 4'b0101;
	mem[2200] = 4'b0101;
	mem[2201] = 4'b0101;
	mem[2202] = 4'b0111;
	mem[2203] = 4'b0110;
	mem[2204] = 4'b0110;
	mem[2205] = 4'b0110;
	mem[2206] = 4'b0110;
	mem[2207] = 4'b0101;
	mem[2208] = 4'b0101;
	mem[2209] = 4'b0110;
	mem[2210] = 4'b0110;
	mem[2211] = 4'b0110;
	mem[2212] = 4'b0110;
	mem[2213] = 4'b1101;
	mem[2214] = 4'b1111;
	mem[2215] = 4'b1111;
	mem[2216] = 4'b1111;
	mem[2217] = 4'b1111;
	mem[2218] = 4'b1111;
	mem[2219] = 4'b1111;
	mem[2220] = 4'b1111;
	mem[2221] = 4'b1111;
	mem[2222] = 4'b1111;
	mem[2223] = 4'b1111;
	mem[2224] = 4'b1111;
	mem[2225] = 4'b1111;
	mem[2226] = 4'b1111;
	mem[2227] = 4'b1111;
	mem[2228] = 4'b1111;
	mem[2229] = 4'b1111;
	mem[2230] = 4'b1010;
	mem[2231] = 4'b0111;
	mem[2232] = 4'b0111;
	mem[2233] = 4'b0111;
	mem[2234] = 4'b0111;
	mem[2235] = 4'b0101;
	mem[2236] = 4'b0011;
	mem[2237] = 4'b0001;
	mem[2238] = 4'b0000;
	mem[2239] = 4'b0000;
	mem[2240] = 4'b0000;
	mem[2241] = 4'b0000;
	mem[2242] = 4'b0000;
	mem[2243] = 4'b0000;
	mem[2244] = 4'b0000;
	mem[2245] = 4'b0000;
	mem[2246] = 4'b0000;
	mem[2247] = 4'b1100;
	mem[2248] = 4'b1111;
	mem[2249] = 4'b1111;
	mem[2250] = 4'b1111;
	mem[2251] = 4'b1111;
	mem[2252] = 4'b1111;
	mem[2253] = 4'b1111;
	mem[2254] = 4'b1111;
	mem[2255] = 4'b1111;
	mem[2256] = 4'b1111;
	mem[2257] = 4'b1111;
	mem[2258] = 4'b1111;
	mem[2259] = 4'b1111;
	mem[2260] = 4'b1111;
	mem[2261] = 4'b1111;
	mem[2262] = 4'b1111;
	mem[2263] = 4'b1110;
	mem[2264] = 4'b0011;
	mem[2265] = 4'b0000;
	mem[2266] = 4'b0000;
	mem[2267] = 4'b0001;
	mem[2268] = 4'b0001;
	mem[2269] = 4'b0000;
	mem[2270] = 4'b0000;
	mem[2271] = 4'b0000;
	mem[2272] = 4'b0000;
	mem[2273] = 4'b0000;
	mem[2274] = 4'b0000;
	mem[2275] = 4'b0000;
	mem[2276] = 4'b0000;
	mem[2277] = 4'b0000;
	mem[2278] = 4'b0000;
	mem[2279] = 4'b0000;
	mem[2280] = 4'b0000;
	mem[2281] = 4'b1010;
	mem[2282] = 4'b1111;
	mem[2283] = 4'b1111;
	mem[2284] = 4'b1111;
	mem[2285] = 4'b1111;
	mem[2286] = 4'b1111;
	mem[2287] = 4'b1111;
	mem[2288] = 4'b1111;
	mem[2289] = 4'b1111;
	mem[2290] = 4'b1111;
	mem[2291] = 4'b1111;
	mem[2292] = 4'b1111;
	mem[2293] = 4'b1111;
	mem[2294] = 4'b1111;
	mem[2295] = 4'b1111;
	mem[2296] = 4'b1111;
	mem[2297] = 4'b1111;
	mem[2298] = 4'b0011;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0111;
	mem[2308] = 4'b1100;
	mem[2309] = 4'b1101;
	mem[2310] = 4'b1101;
	mem[2311] = 4'b1101;
	mem[2312] = 4'b1101;
	mem[2313] = 4'b1101;
	mem[2314] = 4'b1101;
	mem[2315] = 4'b1101;
	mem[2316] = 4'b1101;
	mem[2317] = 4'b1101;
	mem[2318] = 4'b1110;
	mem[2319] = 4'b1110;
	mem[2320] = 4'b1110;
	mem[2321] = 4'b1110;
	mem[2322] = 4'b1110;
	mem[2323] = 4'b1110;
	mem[2324] = 4'b1000;
	mem[2325] = 4'b0110;
	mem[2326] = 4'b0110;
	mem[2327] = 4'b0110;
	mem[2328] = 4'b0101;
	mem[2329] = 4'b0101;
	mem[2330] = 4'b0110;
	mem[2331] = 4'b0110;
	mem[2332] = 4'b0110;
	mem[2333] = 4'b0110;
	mem[2334] = 4'b0110;
	mem[2335] = 4'b0110;
	mem[2336] = 4'b0101;
	mem[2337] = 4'b0110;
	mem[2338] = 4'b0111;
	mem[2339] = 4'b0110;
	mem[2340] = 4'b0110;
	mem[2341] = 4'b1101;
	mem[2342] = 4'b1111;
	mem[2343] = 4'b1111;
	mem[2344] = 4'b1111;
	mem[2345] = 4'b1111;
	mem[2346] = 4'b1111;
	mem[2347] = 4'b1111;
	mem[2348] = 4'b1111;
	mem[2349] = 4'b1111;
	mem[2350] = 4'b1111;
	mem[2351] = 4'b1111;
	mem[2352] = 4'b1111;
	mem[2353] = 4'b1111;
	mem[2354] = 4'b1111;
	mem[2355] = 4'b1111;
	mem[2356] = 4'b1111;
	mem[2357] = 4'b1111;
	mem[2358] = 4'b1010;
	mem[2359] = 4'b0111;
	mem[2360] = 4'b0101;
	mem[2361] = 4'b0011;
	mem[2362] = 4'b0001;
	mem[2363] = 4'b0000;
	mem[2364] = 4'b0000;
	mem[2365] = 4'b0000;
	mem[2366] = 4'b0000;
	mem[2367] = 4'b0000;
	mem[2368] = 4'b0000;
	mem[2369] = 4'b0000;
	mem[2370] = 4'b0000;
	mem[2371] = 4'b0000;
	mem[2372] = 4'b0000;
	mem[2373] = 4'b0000;
	mem[2374] = 4'b0000;
	mem[2375] = 4'b1100;
	mem[2376] = 4'b1111;
	mem[2377] = 4'b1111;
	mem[2378] = 4'b1111;
	mem[2379] = 4'b1111;
	mem[2380] = 4'b1111;
	mem[2381] = 4'b1111;
	mem[2382] = 4'b1111;
	mem[2383] = 4'b1111;
	mem[2384] = 4'b1111;
	mem[2385] = 4'b1111;
	mem[2386] = 4'b1111;
	mem[2387] = 4'b1111;
	mem[2388] = 4'b1111;
	mem[2389] = 4'b1111;
	mem[2390] = 4'b1111;
	mem[2391] = 4'b1111;
	mem[2392] = 4'b0100;
	mem[2393] = 4'b0001;
	mem[2394] = 4'b0001;
	mem[2395] = 4'b0000;
	mem[2396] = 4'b0000;
	mem[2397] = 4'b0000;
	mem[2398] = 4'b0000;
	mem[2399] = 4'b0000;
	mem[2400] = 4'b0000;
	mem[2401] = 4'b0000;
	mem[2402] = 4'b0000;
	mem[2403] = 4'b0000;
	mem[2404] = 4'b0000;
	mem[2405] = 4'b0000;
	mem[2406] = 4'b0000;
	mem[2407] = 4'b0000;
	mem[2408] = 4'b0000;
	mem[2409] = 4'b1010;
	mem[2410] = 4'b1111;
	mem[2411] = 4'b1111;
	mem[2412] = 4'b1111;
	mem[2413] = 4'b1111;
	mem[2414] = 4'b1111;
	mem[2415] = 4'b1111;
	mem[2416] = 4'b1111;
	mem[2417] = 4'b1111;
	mem[2418] = 4'b1111;
	mem[2419] = 4'b1111;
	mem[2420] = 4'b1111;
	mem[2421] = 4'b1111;
	mem[2422] = 4'b1111;
	mem[2423] = 4'b1111;
	mem[2424] = 4'b1111;
	mem[2425] = 4'b1111;
	mem[2426] = 4'b0011;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0111;
	mem[2436] = 4'b1100;
	mem[2437] = 4'b1101;
	mem[2438] = 4'b1101;
	mem[2439] = 4'b1101;
	mem[2440] = 4'b1101;
	mem[2441] = 4'b1101;
	mem[2442] = 4'b1101;
	mem[2443] = 4'b1101;
	mem[2444] = 4'b1110;
	mem[2445] = 4'b1110;
	mem[2446] = 4'b1110;
	mem[2447] = 4'b1110;
	mem[2448] = 4'b1110;
	mem[2449] = 4'b1110;
	mem[2450] = 4'b1110;
	mem[2451] = 4'b1110;
	mem[2452] = 4'b1000;
	mem[2453] = 4'b0110;
	mem[2454] = 4'b0110;
	mem[2455] = 4'b0110;
	mem[2456] = 4'b0110;
	mem[2457] = 4'b0101;
	mem[2458] = 4'b0101;
	mem[2459] = 4'b0110;
	mem[2460] = 4'b0110;
	mem[2461] = 4'b0110;
	mem[2462] = 4'b0110;
	mem[2463] = 4'b0110;
	mem[2464] = 4'b0111;
	mem[2465] = 4'b0111;
	mem[2466] = 4'b0110;
	mem[2467] = 4'b0110;
	mem[2468] = 4'b0110;
	mem[2469] = 4'b1101;
	mem[2470] = 4'b1111;
	mem[2471] = 4'b1111;
	mem[2472] = 4'b1111;
	mem[2473] = 4'b1111;
	mem[2474] = 4'b1111;
	mem[2475] = 4'b1111;
	mem[2476] = 4'b1111;
	mem[2477] = 4'b1111;
	mem[2478] = 4'b1111;
	mem[2479] = 4'b1111;
	mem[2480] = 4'b1111;
	mem[2481] = 4'b1111;
	mem[2482] = 4'b1111;
	mem[2483] = 4'b1111;
	mem[2484] = 4'b1111;
	mem[2485] = 4'b1111;
	mem[2486] = 4'b1000;
	mem[2487] = 4'b0001;
	mem[2488] = 4'b0000;
	mem[2489] = 4'b0000;
	mem[2490] = 4'b0000;
	mem[2491] = 4'b0000;
	mem[2492] = 4'b0000;
	mem[2493] = 4'b0000;
	mem[2494] = 4'b0000;
	mem[2495] = 4'b0000;
	mem[2496] = 4'b0000;
	mem[2497] = 4'b0000;
	mem[2498] = 4'b0000;
	mem[2499] = 4'b0000;
	mem[2500] = 4'b0000;
	mem[2501] = 4'b0000;
	mem[2502] = 4'b0000;
	mem[2503] = 4'b1100;
	mem[2504] = 4'b1111;
	mem[2505] = 4'b1111;
	mem[2506] = 4'b1111;
	mem[2507] = 4'b1111;
	mem[2508] = 4'b1111;
	mem[2509] = 4'b1111;
	mem[2510] = 4'b1111;
	mem[2511] = 4'b1111;
	mem[2512] = 4'b1111;
	mem[2513] = 4'b1111;
	mem[2514] = 4'b1111;
	mem[2515] = 4'b1111;
	mem[2516] = 4'b1110;
	mem[2517] = 4'b1111;
	mem[2518] = 4'b1111;
	mem[2519] = 4'b1111;
	mem[2520] = 4'b0100;
	mem[2521] = 4'b0000;
	mem[2522] = 4'b0000;
	mem[2523] = 4'b0000;
	mem[2524] = 4'b0000;
	mem[2525] = 4'b0000;
	mem[2526] = 4'b0000;
	mem[2527] = 4'b0000;
	mem[2528] = 4'b0000;
	mem[2529] = 4'b0000;
	mem[2530] = 4'b0000;
	mem[2531] = 4'b0000;
	mem[2532] = 4'b0000;
	mem[2533] = 4'b0000;
	mem[2534] = 4'b0000;
	mem[2535] = 4'b0000;
	mem[2536] = 4'b0000;
	mem[2537] = 4'b1010;
	mem[2538] = 4'b1111;
	mem[2539] = 4'b1111;
	mem[2540] = 4'b1111;
	mem[2541] = 4'b1111;
	mem[2542] = 4'b1111;
	mem[2543] = 4'b1111;
	mem[2544] = 4'b1111;
	mem[2545] = 4'b1111;
	mem[2546] = 4'b1111;
	mem[2547] = 4'b1111;
	mem[2548] = 4'b1111;
	mem[2549] = 4'b1111;
	mem[2550] = 4'b1111;
	mem[2551] = 4'b1111;
	mem[2552] = 4'b1111;
	mem[2553] = 4'b1111;
	mem[2554] = 4'b0011;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b0111;
	mem[2564] = 4'b1100;
	mem[2565] = 4'b1101;
	mem[2566] = 4'b1101;
	mem[2567] = 4'b1101;
	mem[2568] = 4'b1101;
	mem[2569] = 4'b1101;
	mem[2570] = 4'b1110;
	mem[2571] = 4'b1110;
	mem[2572] = 4'b1110;
	mem[2573] = 4'b1110;
	mem[2574] = 4'b1110;
	mem[2575] = 4'b1110;
	mem[2576] = 4'b1110;
	mem[2577] = 4'b1110;
	mem[2578] = 4'b1101;
	mem[2579] = 4'b1101;
	mem[2580] = 4'b0111;
	mem[2581] = 4'b0110;
	mem[2582] = 4'b0110;
	mem[2583] = 4'b0110;
	mem[2584] = 4'b0110;
	mem[2585] = 4'b0110;
	mem[2586] = 4'b0101;
	mem[2587] = 4'b0101;
	mem[2588] = 4'b0110;
	mem[2589] = 4'b0110;
	mem[2590] = 4'b0110;
	mem[2591] = 4'b0110;
	mem[2592] = 4'b0110;
	mem[2593] = 4'b0110;
	mem[2594] = 4'b0110;
	mem[2595] = 4'b0110;
	mem[2596] = 4'b0110;
	mem[2597] = 4'b1101;
	mem[2598] = 4'b1111;
	mem[2599] = 4'b1111;
	mem[2600] = 4'b1111;
	mem[2601] = 4'b1111;
	mem[2602] = 4'b1111;
	mem[2603] = 4'b1111;
	mem[2604] = 4'b1111;
	mem[2605] = 4'b1111;
	mem[2606] = 4'b1111;
	mem[2607] = 4'b1111;
	mem[2608] = 4'b1111;
	mem[2609] = 4'b1111;
	mem[2610] = 4'b1111;
	mem[2611] = 4'b1111;
	mem[2612] = 4'b1111;
	mem[2613] = 4'b1111;
	mem[2614] = 4'b0110;
	mem[2615] = 4'b0000;
	mem[2616] = 4'b0000;
	mem[2617] = 4'b0000;
	mem[2618] = 4'b0000;
	mem[2619] = 4'b0000;
	mem[2620] = 4'b0000;
	mem[2621] = 4'b0000;
	mem[2622] = 4'b0000;
	mem[2623] = 4'b0000;
	mem[2624] = 4'b0000;
	mem[2625] = 4'b0000;
	mem[2626] = 4'b0000;
	mem[2627] = 4'b0000;
	mem[2628] = 4'b0000;
	mem[2629] = 4'b0000;
	mem[2630] = 4'b0000;
	mem[2631] = 4'b1011;
	mem[2632] = 4'b1111;
	mem[2633] = 4'b1111;
	mem[2634] = 4'b1111;
	mem[2635] = 4'b1111;
	mem[2636] = 4'b1111;
	mem[2637] = 4'b1111;
	mem[2638] = 4'b1111;
	mem[2639] = 4'b1111;
	mem[2640] = 4'b1111;
	mem[2641] = 4'b1111;
	mem[2642] = 4'b1111;
	mem[2643] = 4'b1111;
	mem[2644] = 4'b1101;
	mem[2645] = 4'b1101;
	mem[2646] = 4'b1111;
	mem[2647] = 4'b1111;
	mem[2648] = 4'b0100;
	mem[2649] = 4'b0000;
	mem[2650] = 4'b0000;
	mem[2651] = 4'b0000;
	mem[2652] = 4'b0000;
	mem[2653] = 4'b0000;
	mem[2654] = 4'b0000;
	mem[2655] = 4'b0000;
	mem[2656] = 4'b0000;
	mem[2657] = 4'b0000;
	mem[2658] = 4'b0000;
	mem[2659] = 4'b0000;
	mem[2660] = 4'b0000;
	mem[2661] = 4'b0000;
	mem[2662] = 4'b0000;
	mem[2663] = 4'b0000;
	mem[2664] = 4'b0000;
	mem[2665] = 4'b1010;
	mem[2666] = 4'b1111;
	mem[2667] = 4'b1111;
	mem[2668] = 4'b1111;
	mem[2669] = 4'b1111;
	mem[2670] = 4'b1111;
	mem[2671] = 4'b1111;
	mem[2672] = 4'b1111;
	mem[2673] = 4'b1111;
	mem[2674] = 4'b1111;
	mem[2675] = 4'b1111;
	mem[2676] = 4'b1111;
	mem[2677] = 4'b1111;
	mem[2678] = 4'b1111;
	mem[2679] = 4'b1111;
	mem[2680] = 4'b1111;
	mem[2681] = 4'b1111;
	mem[2682] = 4'b0011;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b0111;
	mem[2692] = 4'b1100;
	mem[2693] = 4'b1101;
	mem[2694] = 4'b1101;
	mem[2695] = 4'b1101;
	mem[2696] = 4'b1110;
	mem[2697] = 4'b1110;
	mem[2698] = 4'b1110;
	mem[2699] = 4'b1110;
	mem[2700] = 4'b1110;
	mem[2701] = 4'b1110;
	mem[2702] = 4'b1110;
	mem[2703] = 4'b1110;
	mem[2704] = 4'b1110;
	mem[2705] = 4'b1101;
	mem[2706] = 4'b1100;
	mem[2707] = 4'b1100;
	mem[2708] = 4'b0111;
	mem[2709] = 4'b0101;
	mem[2710] = 4'b0101;
	mem[2711] = 4'b0110;
	mem[2712] = 4'b0110;
	mem[2713] = 4'b0110;
	mem[2714] = 4'b0110;
	mem[2715] = 4'b0101;
	mem[2716] = 4'b0101;
	mem[2717] = 4'b0110;
	mem[2718] = 4'b0110;
	mem[2719] = 4'b0110;
	mem[2720] = 4'b0110;
	mem[2721] = 4'b0110;
	mem[2722] = 4'b0110;
	mem[2723] = 4'b0110;
	mem[2724] = 4'b0110;
	mem[2725] = 4'b1101;
	mem[2726] = 4'b1111;
	mem[2727] = 4'b1111;
	mem[2728] = 4'b1111;
	mem[2729] = 4'b1111;
	mem[2730] = 4'b1111;
	mem[2731] = 4'b1111;
	mem[2732] = 4'b1111;
	mem[2733] = 4'b1111;
	mem[2734] = 4'b1111;
	mem[2735] = 4'b1111;
	mem[2736] = 4'b1111;
	mem[2737] = 4'b1111;
	mem[2738] = 4'b1111;
	mem[2739] = 4'b1111;
	mem[2740] = 4'b1111;
	mem[2741] = 4'b1111;
	mem[2742] = 4'b0110;
	mem[2743] = 4'b0000;
	mem[2744] = 4'b0000;
	mem[2745] = 4'b0000;
	mem[2746] = 4'b0000;
	mem[2747] = 4'b0000;
	mem[2748] = 4'b0000;
	mem[2749] = 4'b0000;
	mem[2750] = 4'b0000;
	mem[2751] = 4'b0000;
	mem[2752] = 4'b0000;
	mem[2753] = 4'b0000;
	mem[2754] = 4'b0000;
	mem[2755] = 4'b0000;
	mem[2756] = 4'b0000;
	mem[2757] = 4'b0000;
	mem[2758] = 4'b0000;
	mem[2759] = 4'b1010;
	mem[2760] = 4'b1111;
	mem[2761] = 4'b1111;
	mem[2762] = 4'b1111;
	mem[2763] = 4'b1111;
	mem[2764] = 4'b1111;
	mem[2765] = 4'b1111;
	mem[2766] = 4'b1111;
	mem[2767] = 4'b1111;
	mem[2768] = 4'b1111;
	mem[2769] = 4'b1111;
	mem[2770] = 4'b1111;
	mem[2771] = 4'b1101;
	mem[2772] = 4'b1101;
	mem[2773] = 4'b1101;
	mem[2774] = 4'b1101;
	mem[2775] = 4'b1111;
	mem[2776] = 4'b0100;
	mem[2777] = 4'b0000;
	mem[2778] = 4'b0000;
	mem[2779] = 4'b0000;
	mem[2780] = 4'b0000;
	mem[2781] = 4'b0000;
	mem[2782] = 4'b0000;
	mem[2783] = 4'b0000;
	mem[2784] = 4'b0000;
	mem[2785] = 4'b0000;
	mem[2786] = 4'b0000;
	mem[2787] = 4'b0000;
	mem[2788] = 4'b0000;
	mem[2789] = 4'b0000;
	mem[2790] = 4'b0000;
	mem[2791] = 4'b0000;
	mem[2792] = 4'b0000;
	mem[2793] = 4'b1010;
	mem[2794] = 4'b1111;
	mem[2795] = 4'b1111;
	mem[2796] = 4'b1111;
	mem[2797] = 4'b1111;
	mem[2798] = 4'b1111;
	mem[2799] = 4'b1111;
	mem[2800] = 4'b1111;
	mem[2801] = 4'b1110;
	mem[2802] = 4'b1101;
	mem[2803] = 4'b1111;
	mem[2804] = 4'b1111;
	mem[2805] = 4'b1111;
	mem[2806] = 4'b1111;
	mem[2807] = 4'b1111;
	mem[2808] = 4'b1111;
	mem[2809] = 4'b1111;
	mem[2810] = 4'b0011;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b0111;
	mem[2820] = 4'b1100;
	mem[2821] = 4'b1101;
	mem[2822] = 4'b1101;
	mem[2823] = 4'b1110;
	mem[2824] = 4'b1110;
	mem[2825] = 4'b1110;
	mem[2826] = 4'b1110;
	mem[2827] = 4'b1110;
	mem[2828] = 4'b1110;
	mem[2829] = 4'b1110;
	mem[2830] = 4'b1110;
	mem[2831] = 4'b1110;
	mem[2832] = 4'b1101;
	mem[2833] = 4'b1100;
	mem[2834] = 4'b1100;
	mem[2835] = 4'b1101;
	mem[2836] = 4'b1000;
	mem[2837] = 4'b0110;
	mem[2838] = 4'b0110;
	mem[2839] = 4'b0101;
	mem[2840] = 4'b0110;
	mem[2841] = 4'b0110;
	mem[2842] = 4'b0110;
	mem[2843] = 4'b0110;
	mem[2844] = 4'b0101;
	mem[2845] = 4'b0110;
	mem[2846] = 4'b0111;
	mem[2847] = 4'b0110;
	mem[2848] = 4'b0110;
	mem[2849] = 4'b0110;
	mem[2850] = 4'b0110;
	mem[2851] = 4'b0110;
	mem[2852] = 4'b0110;
	mem[2853] = 4'b1101;
	mem[2854] = 4'b1111;
	mem[2855] = 4'b1111;
	mem[2856] = 4'b1111;
	mem[2857] = 4'b1111;
	mem[2858] = 4'b1111;
	mem[2859] = 4'b1111;
	mem[2860] = 4'b1111;
	mem[2861] = 4'b1111;
	mem[2862] = 4'b1111;
	mem[2863] = 4'b1111;
	mem[2864] = 4'b1111;
	mem[2865] = 4'b1111;
	mem[2866] = 4'b1111;
	mem[2867] = 4'b1111;
	mem[2868] = 4'b1111;
	mem[2869] = 4'b1111;
	mem[2870] = 4'b0110;
	mem[2871] = 4'b0000;
	mem[2872] = 4'b0000;
	mem[2873] = 4'b0000;
	mem[2874] = 4'b0000;
	mem[2875] = 4'b0000;
	mem[2876] = 4'b0000;
	mem[2877] = 4'b0000;
	mem[2878] = 4'b0000;
	mem[2879] = 4'b0000;
	mem[2880] = 4'b0000;
	mem[2881] = 4'b0000;
	mem[2882] = 4'b0000;
	mem[2883] = 4'b0000;
	mem[2884] = 4'b0000;
	mem[2885] = 4'b0000;
	mem[2886] = 4'b0000;
	mem[2887] = 4'b1010;
	mem[2888] = 4'b1101;
	mem[2889] = 4'b1111;
	mem[2890] = 4'b1111;
	mem[2891] = 4'b1111;
	mem[2892] = 4'b1111;
	mem[2893] = 4'b1111;
	mem[2894] = 4'b1111;
	mem[2895] = 4'b1111;
	mem[2896] = 4'b1111;
	mem[2897] = 4'b1111;
	mem[2898] = 4'b1101;
	mem[2899] = 4'b1101;
	mem[2900] = 4'b1101;
	mem[2901] = 4'b1101;
	mem[2902] = 4'b1110;
	mem[2903] = 4'b1111;
	mem[2904] = 4'b0100;
	mem[2905] = 4'b0000;
	mem[2906] = 4'b0000;
	mem[2907] = 4'b0000;
	mem[2908] = 4'b0000;
	mem[2909] = 4'b0000;
	mem[2910] = 4'b0000;
	mem[2911] = 4'b0000;
	mem[2912] = 4'b0000;
	mem[2913] = 4'b0000;
	mem[2914] = 4'b0000;
	mem[2915] = 4'b0000;
	mem[2916] = 4'b0000;
	mem[2917] = 4'b0000;
	mem[2918] = 4'b0000;
	mem[2919] = 4'b0000;
	mem[2920] = 4'b0000;
	mem[2921] = 4'b1010;
	mem[2922] = 4'b1111;
	mem[2923] = 4'b1111;
	mem[2924] = 4'b1111;
	mem[2925] = 4'b1111;
	mem[2926] = 4'b1111;
	mem[2927] = 4'b1111;
	mem[2928] = 4'b1111;
	mem[2929] = 4'b1110;
	mem[2930] = 4'b1101;
	mem[2931] = 4'b1101;
	mem[2932] = 4'b1111;
	mem[2933] = 4'b1111;
	mem[2934] = 4'b1111;
	mem[2935] = 4'b1111;
	mem[2936] = 4'b1111;
	mem[2937] = 4'b1111;
	mem[2938] = 4'b0011;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b0111;
	mem[2948] = 4'b1100;
	mem[2949] = 4'b1101;
	mem[2950] = 4'b1110;
	mem[2951] = 4'b1110;
	mem[2952] = 4'b1110;
	mem[2953] = 4'b1110;
	mem[2954] = 4'b1110;
	mem[2955] = 4'b1110;
	mem[2956] = 4'b1110;
	mem[2957] = 4'b1110;
	mem[2958] = 4'b1110;
	mem[2959] = 4'b1110;
	mem[2960] = 4'b1101;
	mem[2961] = 4'b1100;
	mem[2962] = 4'b1100;
	mem[2963] = 4'b1110;
	mem[2964] = 4'b1000;
	mem[2965] = 4'b0110;
	mem[2966] = 4'b0110;
	mem[2967] = 4'b0110;
	mem[2968] = 4'b0101;
	mem[2969] = 4'b0111;
	mem[2970] = 4'b0110;
	mem[2971] = 4'b0110;
	mem[2972] = 4'b0111;
	mem[2973] = 4'b0111;
	mem[2974] = 4'b0111;
	mem[2975] = 4'b0110;
	mem[2976] = 4'b0110;
	mem[2977] = 4'b0110;
	mem[2978] = 4'b0110;
	mem[2979] = 4'b0110;
	mem[2980] = 4'b0110;
	mem[2981] = 4'b1101;
	mem[2982] = 4'b1111;
	mem[2983] = 4'b1111;
	mem[2984] = 4'b1111;
	mem[2985] = 4'b1111;
	mem[2986] = 4'b1111;
	mem[2987] = 4'b1111;
	mem[2988] = 4'b1111;
	mem[2989] = 4'b1111;
	mem[2990] = 4'b1111;
	mem[2991] = 4'b1111;
	mem[2992] = 4'b1111;
	mem[2993] = 4'b1111;
	mem[2994] = 4'b1111;
	mem[2995] = 4'b1111;
	mem[2996] = 4'b1111;
	mem[2997] = 4'b1111;
	mem[2998] = 4'b0110;
	mem[2999] = 4'b0000;
	mem[3000] = 4'b0000;
	mem[3001] = 4'b0000;
	mem[3002] = 4'b0000;
	mem[3003] = 4'b0000;
	mem[3004] = 4'b0000;
	mem[3005] = 4'b0000;
	mem[3006] = 4'b0000;
	mem[3007] = 4'b0000;
	mem[3008] = 4'b0000;
	mem[3009] = 4'b0000;
	mem[3010] = 4'b0000;
	mem[3011] = 4'b0000;
	mem[3012] = 4'b0000;
	mem[3013] = 4'b0000;
	mem[3014] = 4'b0000;
	mem[3015] = 4'b1010;
	mem[3016] = 4'b1101;
	mem[3017] = 4'b1101;
	mem[3018] = 4'b1111;
	mem[3019] = 4'b1111;
	mem[3020] = 4'b1111;
	mem[3021] = 4'b1111;
	mem[3022] = 4'b1111;
	mem[3023] = 4'b1111;
	mem[3024] = 4'b1111;
	mem[3025] = 4'b1101;
	mem[3026] = 4'b1101;
	mem[3027] = 4'b1101;
	mem[3028] = 4'b1101;
	mem[3029] = 4'b1110;
	mem[3030] = 4'b1111;
	mem[3031] = 4'b1111;
	mem[3032] = 4'b0100;
	mem[3033] = 4'b0000;
	mem[3034] = 4'b0000;
	mem[3035] = 4'b0000;
	mem[3036] = 4'b0000;
	mem[3037] = 4'b0000;
	mem[3038] = 4'b0000;
	mem[3039] = 4'b0000;
	mem[3040] = 4'b0000;
	mem[3041] = 4'b0000;
	mem[3042] = 4'b0000;
	mem[3043] = 4'b0000;
	mem[3044] = 4'b0000;
	mem[3045] = 4'b0000;
	mem[3046] = 4'b0000;
	mem[3047] = 4'b0000;
	mem[3048] = 4'b0000;
	mem[3049] = 4'b1010;
	mem[3050] = 4'b1111;
	mem[3051] = 4'b1111;
	mem[3052] = 4'b1111;
	mem[3053] = 4'b1111;
	mem[3054] = 4'b1111;
	mem[3055] = 4'b1111;
	mem[3056] = 4'b1111;
	mem[3057] = 4'b1111;
	mem[3058] = 4'b1110;
	mem[3059] = 4'b1101;
	mem[3060] = 4'b1101;
	mem[3061] = 4'b1111;
	mem[3062] = 4'b1111;
	mem[3063] = 4'b1111;
	mem[3064] = 4'b1111;
	mem[3065] = 4'b1111;
	mem[3066] = 4'b0011;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b0111;
	mem[3076] = 4'b1100;
	mem[3077] = 4'b1101;
	mem[3078] = 4'b1110;
	mem[3079] = 4'b1110;
	mem[3080] = 4'b1110;
	mem[3081] = 4'b1110;
	mem[3082] = 4'b1110;
	mem[3083] = 4'b1110;
	mem[3084] = 4'b1110;
	mem[3085] = 4'b1110;
	mem[3086] = 4'b1110;
	mem[3087] = 4'b1110;
	mem[3088] = 4'b1101;
	mem[3089] = 4'b1100;
	mem[3090] = 4'b1101;
	mem[3091] = 4'b1110;
	mem[3092] = 4'b1000;
	mem[3093] = 4'b0110;
	mem[3094] = 4'b0110;
	mem[3095] = 4'b0110;
	mem[3096] = 4'b0101;
	mem[3097] = 4'b0110;
	mem[3098] = 4'b0111;
	mem[3099] = 4'b0110;
	mem[3100] = 4'b0110;
	mem[3101] = 4'b0110;
	mem[3102] = 4'b0110;
	mem[3103] = 4'b0110;
	mem[3104] = 4'b0110;
	mem[3105] = 4'b0110;
	mem[3106] = 4'b0110;
	mem[3107] = 4'b0110;
	mem[3108] = 4'b0110;
	mem[3109] = 4'b1101;
	mem[3110] = 4'b1111;
	mem[3111] = 4'b1111;
	mem[3112] = 4'b1111;
	mem[3113] = 4'b1111;
	mem[3114] = 4'b1111;
	mem[3115] = 4'b1111;
	mem[3116] = 4'b1111;
	mem[3117] = 4'b1111;
	mem[3118] = 4'b1111;
	mem[3119] = 4'b1111;
	mem[3120] = 4'b1111;
	mem[3121] = 4'b1111;
	mem[3122] = 4'b1111;
	mem[3123] = 4'b1111;
	mem[3124] = 4'b1111;
	mem[3125] = 4'b1111;
	mem[3126] = 4'b0110;
	mem[3127] = 4'b0000;
	mem[3128] = 4'b0000;
	mem[3129] = 4'b0000;
	mem[3130] = 4'b0000;
	mem[3131] = 4'b0000;
	mem[3132] = 4'b0000;
	mem[3133] = 4'b0000;
	mem[3134] = 4'b0000;
	mem[3135] = 4'b0000;
	mem[3136] = 4'b0000;
	mem[3137] = 4'b0000;
	mem[3138] = 4'b0000;
	mem[3139] = 4'b0000;
	mem[3140] = 4'b0000;
	mem[3141] = 4'b0000;
	mem[3142] = 4'b0000;
	mem[3143] = 4'b1010;
	mem[3144] = 4'b1101;
	mem[3145] = 4'b1101;
	mem[3146] = 4'b1101;
	mem[3147] = 4'b1111;
	mem[3148] = 4'b1111;
	mem[3149] = 4'b1111;
	mem[3150] = 4'b1111;
	mem[3151] = 4'b1111;
	mem[3152] = 4'b1101;
	mem[3153] = 4'b1101;
	mem[3154] = 4'b1101;
	mem[3155] = 4'b1101;
	mem[3156] = 4'b1110;
	mem[3157] = 4'b1111;
	mem[3158] = 4'b1111;
	mem[3159] = 4'b1111;
	mem[3160] = 4'b0100;
	mem[3161] = 4'b0000;
	mem[3162] = 4'b0000;
	mem[3163] = 4'b0000;
	mem[3164] = 4'b0000;
	mem[3165] = 4'b0000;
	mem[3166] = 4'b0000;
	mem[3167] = 4'b0000;
	mem[3168] = 4'b0000;
	mem[3169] = 4'b0000;
	mem[3170] = 4'b0000;
	mem[3171] = 4'b0000;
	mem[3172] = 4'b0000;
	mem[3173] = 4'b0000;
	mem[3174] = 4'b0000;
	mem[3175] = 4'b0000;
	mem[3176] = 4'b0000;
	mem[3177] = 4'b1010;
	mem[3178] = 4'b1111;
	mem[3179] = 4'b1111;
	mem[3180] = 4'b1111;
	mem[3181] = 4'b1111;
	mem[3182] = 4'b1111;
	mem[3183] = 4'b1111;
	mem[3184] = 4'b1111;
	mem[3185] = 4'b1111;
	mem[3186] = 4'b1111;
	mem[3187] = 4'b1110;
	mem[3188] = 4'b1101;
	mem[3189] = 4'b1101;
	mem[3190] = 4'b1111;
	mem[3191] = 4'b1111;
	mem[3192] = 4'b1111;
	mem[3193] = 4'b1111;
	mem[3194] = 4'b0011;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b0111;
	mem[3204] = 4'b1100;
	mem[3205] = 4'b1101;
	mem[3206] = 4'b1110;
	mem[3207] = 4'b1110;
	mem[3208] = 4'b1110;
	mem[3209] = 4'b1110;
	mem[3210] = 4'b1110;
	mem[3211] = 4'b1110;
	mem[3212] = 4'b1110;
	mem[3213] = 4'b1110;
	mem[3214] = 4'b1110;
	mem[3215] = 4'b1110;
	mem[3216] = 4'b1101;
	mem[3217] = 4'b1100;
	mem[3218] = 4'b1100;
	mem[3219] = 4'b1110;
	mem[3220] = 4'b1000;
	mem[3221] = 4'b0110;
	mem[3222] = 4'b0110;
	mem[3223] = 4'b0110;
	mem[3224] = 4'b0101;
	mem[3225] = 4'b0110;
	mem[3226] = 4'b0111;
	mem[3227] = 4'b0110;
	mem[3228] = 4'b0110;
	mem[3229] = 4'b0110;
	mem[3230] = 4'b0110;
	mem[3231] = 4'b0110;
	mem[3232] = 4'b0110;
	mem[3233] = 4'b0110;
	mem[3234] = 4'b0110;
	mem[3235] = 4'b0110;
	mem[3236] = 4'b0110;
	mem[3237] = 4'b1101;
	mem[3238] = 4'b1111;
	mem[3239] = 4'b1111;
	mem[3240] = 4'b1111;
	mem[3241] = 4'b1111;
	mem[3242] = 4'b1111;
	mem[3243] = 4'b1111;
	mem[3244] = 4'b1111;
	mem[3245] = 4'b1111;
	mem[3246] = 4'b1111;
	mem[3247] = 4'b1111;
	mem[3248] = 4'b1111;
	mem[3249] = 4'b1111;
	mem[3250] = 4'b1111;
	mem[3251] = 4'b1111;
	mem[3252] = 4'b1111;
	mem[3253] = 4'b1111;
	mem[3254] = 4'b0110;
	mem[3255] = 4'b0000;
	mem[3256] = 4'b0000;
	mem[3257] = 4'b0000;
	mem[3258] = 4'b0000;
	mem[3259] = 4'b0000;
	mem[3260] = 4'b0000;
	mem[3261] = 4'b0000;
	mem[3262] = 4'b0000;
	mem[3263] = 4'b0000;
	mem[3264] = 4'b0000;
	mem[3265] = 4'b0000;
	mem[3266] = 4'b0000;
	mem[3267] = 4'b0000;
	mem[3268] = 4'b0000;
	mem[3269] = 4'b0000;
	mem[3270] = 4'b0000;
	mem[3271] = 4'b1010;
	mem[3272] = 4'b1101;
	mem[3273] = 4'b1101;
	mem[3274] = 4'b1101;
	mem[3275] = 4'b1101;
	mem[3276] = 4'b1111;
	mem[3277] = 4'b1111;
	mem[3278] = 4'b1111;
	mem[3279] = 4'b1101;
	mem[3280] = 4'b1101;
	mem[3281] = 4'b1101;
	mem[3282] = 4'b1101;
	mem[3283] = 4'b1110;
	mem[3284] = 4'b1111;
	mem[3285] = 4'b1111;
	mem[3286] = 4'b1111;
	mem[3287] = 4'b1111;
	mem[3288] = 4'b0100;
	mem[3289] = 4'b0000;
	mem[3290] = 4'b0000;
	mem[3291] = 4'b0000;
	mem[3292] = 4'b0000;
	mem[3293] = 4'b0000;
	mem[3294] = 4'b0000;
	mem[3295] = 4'b0000;
	mem[3296] = 4'b0000;
	mem[3297] = 4'b0000;
	mem[3298] = 4'b0000;
	mem[3299] = 4'b0000;
	mem[3300] = 4'b0000;
	mem[3301] = 4'b0000;
	mem[3302] = 4'b0000;
	mem[3303] = 4'b0000;
	mem[3304] = 4'b0000;
	mem[3305] = 4'b1010;
	mem[3306] = 4'b1111;
	mem[3307] = 4'b1111;
	mem[3308] = 4'b1111;
	mem[3309] = 4'b1111;
	mem[3310] = 4'b1111;
	mem[3311] = 4'b1111;
	mem[3312] = 4'b1111;
	mem[3313] = 4'b1111;
	mem[3314] = 4'b1110;
	mem[3315] = 4'b1110;
	mem[3316] = 4'b1101;
	mem[3317] = 4'b1101;
	mem[3318] = 4'b1101;
	mem[3319] = 4'b1111;
	mem[3320] = 4'b1111;
	mem[3321] = 4'b1111;
	mem[3322] = 4'b0011;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b0111;
	mem[3332] = 4'b1100;
	mem[3333] = 4'b1101;
	mem[3334] = 4'b1110;
	mem[3335] = 4'b1110;
	mem[3336] = 4'b1110;
	mem[3337] = 4'b1110;
	mem[3338] = 4'b1110;
	mem[3339] = 4'b1110;
	mem[3340] = 4'b1110;
	mem[3341] = 4'b1101;
	mem[3342] = 4'b1110;
	mem[3343] = 4'b1110;
	mem[3344] = 4'b1101;
	mem[3345] = 4'b1100;
	mem[3346] = 4'b1100;
	mem[3347] = 4'b1100;
	mem[3348] = 4'b1000;
	mem[3349] = 4'b0110;
	mem[3350] = 4'b0110;
	mem[3351] = 4'b0110;
	mem[3352] = 4'b0110;
	mem[3353] = 4'b0111;
	mem[3354] = 4'b0111;
	mem[3355] = 4'b0110;
	mem[3356] = 4'b0110;
	mem[3357] = 4'b0110;
	mem[3358] = 4'b0110;
	mem[3359] = 4'b0110;
	mem[3360] = 4'b0110;
	mem[3361] = 4'b0110;
	mem[3362] = 4'b0110;
	mem[3363] = 4'b0110;
	mem[3364] = 4'b0110;
	mem[3365] = 4'b1101;
	mem[3366] = 4'b1111;
	mem[3367] = 4'b1111;
	mem[3368] = 4'b1111;
	mem[3369] = 4'b1111;
	mem[3370] = 4'b1111;
	mem[3371] = 4'b1111;
	mem[3372] = 4'b1111;
	mem[3373] = 4'b1111;
	mem[3374] = 4'b1111;
	mem[3375] = 4'b1111;
	mem[3376] = 4'b1111;
	mem[3377] = 4'b1111;
	mem[3378] = 4'b1111;
	mem[3379] = 4'b1111;
	mem[3380] = 4'b1111;
	mem[3381] = 4'b1111;
	mem[3382] = 4'b0110;
	mem[3383] = 4'b0000;
	mem[3384] = 4'b0000;
	mem[3385] = 4'b0000;
	mem[3386] = 4'b0000;
	mem[3387] = 4'b0000;
	mem[3388] = 4'b0000;
	mem[3389] = 4'b0000;
	mem[3390] = 4'b0000;
	mem[3391] = 4'b0000;
	mem[3392] = 4'b0000;
	mem[3393] = 4'b0000;
	mem[3394] = 4'b0000;
	mem[3395] = 4'b0000;
	mem[3396] = 4'b0000;
	mem[3397] = 4'b0000;
	mem[3398] = 4'b0000;
	mem[3399] = 4'b1011;
	mem[3400] = 4'b1101;
	mem[3401] = 4'b1101;
	mem[3402] = 4'b1101;
	mem[3403] = 4'b1101;
	mem[3404] = 4'b1101;
	mem[3405] = 4'b1110;
	mem[3406] = 4'b1101;
	mem[3407] = 4'b1101;
	mem[3408] = 4'b1101;
	mem[3409] = 4'b1101;
	mem[3410] = 4'b1110;
	mem[3411] = 4'b1111;
	mem[3412] = 4'b1111;
	mem[3413] = 4'b1111;
	mem[3414] = 4'b1111;
	mem[3415] = 4'b1111;
	mem[3416] = 4'b0100;
	mem[3417] = 4'b0000;
	mem[3418] = 4'b0000;
	mem[3419] = 4'b0000;
	mem[3420] = 4'b0000;
	mem[3421] = 4'b0000;
	mem[3422] = 4'b0000;
	mem[3423] = 4'b0000;
	mem[3424] = 4'b0000;
	mem[3425] = 4'b0000;
	mem[3426] = 4'b0000;
	mem[3427] = 4'b0000;
	mem[3428] = 4'b0000;
	mem[3429] = 4'b0000;
	mem[3430] = 4'b0000;
	mem[3431] = 4'b0000;
	mem[3432] = 4'b0000;
	mem[3433] = 4'b1010;
	mem[3434] = 4'b1111;
	mem[3435] = 4'b1111;
	mem[3436] = 4'b1111;
	mem[3437] = 4'b1111;
	mem[3438] = 4'b1111;
	mem[3439] = 4'b1111;
	mem[3440] = 4'b1111;
	mem[3441] = 4'b1110;
	mem[3442] = 4'b1101;
	mem[3443] = 4'b1110;
	mem[3444] = 4'b1111;
	mem[3445] = 4'b1110;
	mem[3446] = 4'b1101;
	mem[3447] = 4'b1101;
	mem[3448] = 4'b1111;
	mem[3449] = 4'b1111;
	mem[3450] = 4'b0011;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b0111;
	mem[3460] = 4'b1100;
	mem[3461] = 4'b1101;
	mem[3462] = 4'b1110;
	mem[3463] = 4'b1110;
	mem[3464] = 4'b1110;
	mem[3465] = 4'b1110;
	mem[3466] = 4'b1110;
	mem[3467] = 4'b1101;
	mem[3468] = 4'b1100;
	mem[3469] = 4'b1100;
	mem[3470] = 4'b1100;
	mem[3471] = 4'b1101;
	mem[3472] = 4'b1110;
	mem[3473] = 4'b1101;
	mem[3474] = 4'b1100;
	mem[3475] = 4'b1100;
	mem[3476] = 4'b0111;
	mem[3477] = 4'b0110;
	mem[3478] = 4'b0110;
	mem[3479] = 4'b0110;
	mem[3480] = 4'b0110;
	mem[3481] = 4'b0111;
	mem[3482] = 4'b0110;
	mem[3483] = 4'b0110;
	mem[3484] = 4'b0110;
	mem[3485] = 4'b0110;
	mem[3486] = 4'b0110;
	mem[3487] = 4'b0110;
	mem[3488] = 4'b0110;
	mem[3489] = 4'b0110;
	mem[3490] = 4'b0110;
	mem[3491] = 4'b0011;
	mem[3492] = 4'b0000;
	mem[3493] = 4'b1100;
	mem[3494] = 4'b1111;
	mem[3495] = 4'b1111;
	mem[3496] = 4'b1111;
	mem[3497] = 4'b1111;
	mem[3498] = 4'b1111;
	mem[3499] = 4'b1111;
	mem[3500] = 4'b1111;
	mem[3501] = 4'b1111;
	mem[3502] = 4'b1111;
	mem[3503] = 4'b1111;
	mem[3504] = 4'b1111;
	mem[3505] = 4'b1111;
	mem[3506] = 4'b1111;
	mem[3507] = 4'b1111;
	mem[3508] = 4'b1111;
	mem[3509] = 4'b1111;
	mem[3510] = 4'b0110;
	mem[3511] = 4'b0000;
	mem[3512] = 4'b0000;
	mem[3513] = 4'b0000;
	mem[3514] = 4'b0000;
	mem[3515] = 4'b0000;
	mem[3516] = 4'b0000;
	mem[3517] = 4'b0000;
	mem[3518] = 4'b0000;
	mem[3519] = 4'b0000;
	mem[3520] = 4'b0000;
	mem[3521] = 4'b0000;
	mem[3522] = 4'b0000;
	mem[3523] = 4'b0000;
	mem[3524] = 4'b0000;
	mem[3525] = 4'b0000;
	mem[3526] = 4'b0000;
	mem[3527] = 4'b1100;
	mem[3528] = 4'b1111;
	mem[3529] = 4'b1101;
	mem[3530] = 4'b1101;
	mem[3531] = 4'b1101;
	mem[3532] = 4'b1101;
	mem[3533] = 4'b1101;
	mem[3534] = 4'b1101;
	mem[3535] = 4'b1101;
	mem[3536] = 4'b1101;
	mem[3537] = 4'b1110;
	mem[3538] = 4'b1111;
	mem[3539] = 4'b1111;
	mem[3540] = 4'b1111;
	mem[3541] = 4'b1111;
	mem[3542] = 4'b1111;
	mem[3543] = 4'b1111;
	mem[3544] = 4'b0100;
	mem[3545] = 4'b0000;
	mem[3546] = 4'b0000;
	mem[3547] = 4'b0000;
	mem[3548] = 4'b0000;
	mem[3549] = 4'b0000;
	mem[3550] = 4'b0000;
	mem[3551] = 4'b0000;
	mem[3552] = 4'b0000;
	mem[3553] = 4'b0000;
	mem[3554] = 4'b0000;
	mem[3555] = 4'b0000;
	mem[3556] = 4'b0000;
	mem[3557] = 4'b0000;
	mem[3558] = 4'b0000;
	mem[3559] = 4'b0000;
	mem[3560] = 4'b0000;
	mem[3561] = 4'b1010;
	mem[3562] = 4'b1111;
	mem[3563] = 4'b1111;
	mem[3564] = 4'b1111;
	mem[3565] = 4'b1111;
	mem[3566] = 4'b1111;
	mem[3567] = 4'b1111;
	mem[3568] = 4'b1110;
	mem[3569] = 4'b1101;
	mem[3570] = 4'b1110;
	mem[3571] = 4'b1111;
	mem[3572] = 4'b1111;
	mem[3573] = 4'b1111;
	mem[3574] = 4'b1110;
	mem[3575] = 4'b1101;
	mem[3576] = 4'b1101;
	mem[3577] = 4'b1110;
	mem[3578] = 4'b0011;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b0111;
	mem[3588] = 4'b1100;
	mem[3589] = 4'b1101;
	mem[3590] = 4'b1110;
	mem[3591] = 4'b1110;
	mem[3592] = 4'b1110;
	mem[3593] = 4'b1110;
	mem[3594] = 4'b1101;
	mem[3595] = 4'b1100;
	mem[3596] = 4'b1100;
	mem[3597] = 4'b1100;
	mem[3598] = 4'b1100;
	mem[3599] = 4'b1110;
	mem[3600] = 4'b1110;
	mem[3601] = 4'b1110;
	mem[3602] = 4'b1101;
	mem[3603] = 4'b1100;
	mem[3604] = 4'b0111;
	mem[3605] = 4'b0110;
	mem[3606] = 4'b0110;
	mem[3607] = 4'b0111;
	mem[3608] = 4'b0111;
	mem[3609] = 4'b0111;
	mem[3610] = 4'b0110;
	mem[3611] = 4'b0110;
	mem[3612] = 4'b0110;
	mem[3613] = 4'b0110;
	mem[3614] = 4'b0110;
	mem[3615] = 4'b0110;
	mem[3616] = 4'b0110;
	mem[3617] = 4'b0010;
	mem[3618] = 4'b0000;
	mem[3619] = 4'b0000;
	mem[3620] = 4'b0000;
	mem[3621] = 4'b1100;
	mem[3622] = 4'b1111;
	mem[3623] = 4'b1111;
	mem[3624] = 4'b1111;
	mem[3625] = 4'b1111;
	mem[3626] = 4'b1111;
	mem[3627] = 4'b1111;
	mem[3628] = 4'b1111;
	mem[3629] = 4'b1111;
	mem[3630] = 4'b1111;
	mem[3631] = 4'b1111;
	mem[3632] = 4'b1111;
	mem[3633] = 4'b1111;
	mem[3634] = 4'b1111;
	mem[3635] = 4'b1111;
	mem[3636] = 4'b1111;
	mem[3637] = 4'b1111;
	mem[3638] = 4'b0110;
	mem[3639] = 4'b0000;
	mem[3640] = 4'b0000;
	mem[3641] = 4'b0000;
	mem[3642] = 4'b0000;
	mem[3643] = 4'b0000;
	mem[3644] = 4'b0000;
	mem[3645] = 4'b0000;
	mem[3646] = 4'b0000;
	mem[3647] = 4'b0000;
	mem[3648] = 4'b0000;
	mem[3649] = 4'b0000;
	mem[3650] = 4'b0000;
	mem[3651] = 4'b0000;
	mem[3652] = 4'b0000;
	mem[3653] = 4'b0000;
	mem[3654] = 4'b0000;
	mem[3655] = 4'b1100;
	mem[3656] = 4'b1111;
	mem[3657] = 4'b1111;
	mem[3658] = 4'b1101;
	mem[3659] = 4'b1101;
	mem[3660] = 4'b1101;
	mem[3661] = 4'b1101;
	mem[3662] = 4'b1101;
	mem[3663] = 4'b1101;
	mem[3664] = 4'b1110;
	mem[3665] = 4'b1111;
	mem[3666] = 4'b1111;
	mem[3667] = 4'b1111;
	mem[3668] = 4'b1111;
	mem[3669] = 4'b1111;
	mem[3670] = 4'b1111;
	mem[3671] = 4'b1111;
	mem[3672] = 4'b0100;
	mem[3673] = 4'b0000;
	mem[3674] = 4'b0000;
	mem[3675] = 4'b0000;
	mem[3676] = 4'b0000;
	mem[3677] = 4'b0000;
	mem[3678] = 4'b0000;
	mem[3679] = 4'b0000;
	mem[3680] = 4'b0000;
	mem[3681] = 4'b0000;
	mem[3682] = 4'b0000;
	mem[3683] = 4'b0000;
	mem[3684] = 4'b0000;
	mem[3685] = 4'b0000;
	mem[3686] = 4'b0000;
	mem[3687] = 4'b0000;
	mem[3688] = 4'b0000;
	mem[3689] = 4'b1010;
	mem[3690] = 4'b1111;
	mem[3691] = 4'b1111;
	mem[3692] = 4'b1111;
	mem[3693] = 4'b1111;
	mem[3694] = 4'b1111;
	mem[3695] = 4'b1111;
	mem[3696] = 4'b1110;
	mem[3697] = 4'b1101;
	mem[3698] = 4'b1111;
	mem[3699] = 4'b1111;
	mem[3700] = 4'b1111;
	mem[3701] = 4'b1111;
	mem[3702] = 4'b1111;
	mem[3703] = 4'b1110;
	mem[3704] = 4'b1101;
	mem[3705] = 4'b1101;
	mem[3706] = 4'b0100;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b0111;
	mem[3716] = 4'b1100;
	mem[3717] = 4'b1101;
	mem[3718] = 4'b1110;
	mem[3719] = 4'b1110;
	mem[3720] = 4'b1110;
	mem[3721] = 4'b1101;
	mem[3722] = 4'b1100;
	mem[3723] = 4'b1100;
	mem[3724] = 4'b1101;
	mem[3725] = 4'b1110;
	mem[3726] = 4'b1110;
	mem[3727] = 4'b1110;
	mem[3728] = 4'b1110;
	mem[3729] = 4'b1101;
	mem[3730] = 4'b1110;
	mem[3731] = 4'b1110;
	mem[3732] = 4'b1000;
	mem[3733] = 4'b0111;
	mem[3734] = 4'b0111;
	mem[3735] = 4'b0111;
	mem[3736] = 4'b0111;
	mem[3737] = 4'b0110;
	mem[3738] = 4'b0110;
	mem[3739] = 4'b0110;
	mem[3740] = 4'b0110;
	mem[3741] = 4'b0110;
	mem[3742] = 4'b0110;
	mem[3743] = 4'b0011;
	mem[3744] = 4'b0000;
	mem[3745] = 4'b0000;
	mem[3746] = 4'b0000;
	mem[3747] = 4'b0000;
	mem[3748] = 4'b0000;
	mem[3749] = 4'b1100;
	mem[3750] = 4'b1111;
	mem[3751] = 4'b1111;
	mem[3752] = 4'b1111;
	mem[3753] = 4'b1111;
	mem[3754] = 4'b1111;
	mem[3755] = 4'b1111;
	mem[3756] = 4'b1111;
	mem[3757] = 4'b1111;
	mem[3758] = 4'b1111;
	mem[3759] = 4'b1111;
	mem[3760] = 4'b1111;
	mem[3761] = 4'b1111;
	mem[3762] = 4'b1111;
	mem[3763] = 4'b1111;
	mem[3764] = 4'b1111;
	mem[3765] = 4'b1111;
	mem[3766] = 4'b0110;
	mem[3767] = 4'b0000;
	mem[3768] = 4'b0000;
	mem[3769] = 4'b0000;
	mem[3770] = 4'b0000;
	mem[3771] = 4'b0000;
	mem[3772] = 4'b0000;
	mem[3773] = 4'b0000;
	mem[3774] = 4'b0000;
	mem[3775] = 4'b0000;
	mem[3776] = 4'b0000;
	mem[3777] = 4'b0000;
	mem[3778] = 4'b0000;
	mem[3779] = 4'b0000;
	mem[3780] = 4'b0000;
	mem[3781] = 4'b0000;
	mem[3782] = 4'b0000;
	mem[3783] = 4'b1100;
	mem[3784] = 4'b1111;
	mem[3785] = 4'b1111;
	mem[3786] = 4'b1111;
	mem[3787] = 4'b1101;
	mem[3788] = 4'b1101;
	mem[3789] = 4'b1101;
	mem[3790] = 4'b1101;
	mem[3791] = 4'b1110;
	mem[3792] = 4'b1111;
	mem[3793] = 4'b1111;
	mem[3794] = 4'b1111;
	mem[3795] = 4'b1111;
	mem[3796] = 4'b1111;
	mem[3797] = 4'b1111;
	mem[3798] = 4'b1111;
	mem[3799] = 4'b1111;
	mem[3800] = 4'b0100;
	mem[3801] = 4'b0000;
	mem[3802] = 4'b0000;
	mem[3803] = 4'b0000;
	mem[3804] = 4'b0000;
	mem[3805] = 4'b0000;
	mem[3806] = 4'b0000;
	mem[3807] = 4'b0000;
	mem[3808] = 4'b0000;
	mem[3809] = 4'b0000;
	mem[3810] = 4'b0000;
	mem[3811] = 4'b0000;
	mem[3812] = 4'b0000;
	mem[3813] = 4'b0000;
	mem[3814] = 4'b0000;
	mem[3815] = 4'b0000;
	mem[3816] = 4'b0000;
	mem[3817] = 4'b1010;
	mem[3818] = 4'b1111;
	mem[3819] = 4'b1111;
	mem[3820] = 4'b1111;
	mem[3821] = 4'b1111;
	mem[3822] = 4'b1111;
	mem[3823] = 4'b1111;
	mem[3824] = 4'b1110;
	mem[3825] = 4'b1101;
	mem[3826] = 4'b1110;
	mem[3827] = 4'b1111;
	mem[3828] = 4'b1111;
	mem[3829] = 4'b1111;
	mem[3830] = 4'b1111;
	mem[3831] = 4'b1110;
	mem[3832] = 4'b1101;
	mem[3833] = 4'b1101;
	mem[3834] = 4'b0100;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b0111;
	mem[3844] = 4'b1100;
	mem[3845] = 4'b1101;
	mem[3846] = 4'b1110;
	mem[3847] = 4'b1110;
	mem[3848] = 4'b1110;
	mem[3849] = 4'b1101;
	mem[3850] = 4'b1100;
	mem[3851] = 4'b1100;
	mem[3852] = 4'b1110;
	mem[3853] = 4'b1110;
	mem[3854] = 4'b1110;
	mem[3855] = 4'b1110;
	mem[3856] = 4'b1101;
	mem[3857] = 4'b1100;
	mem[3858] = 4'b1101;
	mem[3859] = 4'b1110;
	mem[3860] = 4'b1000;
	mem[3861] = 4'b0110;
	mem[3862] = 4'b0111;
	mem[3863] = 4'b0110;
	mem[3864] = 4'b0110;
	mem[3865] = 4'b0110;
	mem[3866] = 4'b0110;
	mem[3867] = 4'b0110;
	mem[3868] = 4'b0110;
	mem[3869] = 4'b0011;
	mem[3870] = 4'b0000;
	mem[3871] = 4'b0000;
	mem[3872] = 4'b0000;
	mem[3873] = 4'b0000;
	mem[3874] = 4'b0000;
	mem[3875] = 4'b0000;
	mem[3876] = 4'b0000;
	mem[3877] = 4'b1100;
	mem[3878] = 4'b1111;
	mem[3879] = 4'b1111;
	mem[3880] = 4'b1111;
	mem[3881] = 4'b1111;
	mem[3882] = 4'b1111;
	mem[3883] = 4'b1111;
	mem[3884] = 4'b1111;
	mem[3885] = 4'b1111;
	mem[3886] = 4'b1111;
	mem[3887] = 4'b1111;
	mem[3888] = 4'b1111;
	mem[3889] = 4'b1111;
	mem[3890] = 4'b1111;
	mem[3891] = 4'b1111;
	mem[3892] = 4'b1111;
	mem[3893] = 4'b1111;
	mem[3894] = 4'b0110;
	mem[3895] = 4'b0000;
	mem[3896] = 4'b0000;
	mem[3897] = 4'b0000;
	mem[3898] = 4'b0000;
	mem[3899] = 4'b0000;
	mem[3900] = 4'b0000;
	mem[3901] = 4'b0000;
	mem[3902] = 4'b0000;
	mem[3903] = 4'b0000;
	mem[3904] = 4'b0000;
	mem[3905] = 4'b0000;
	mem[3906] = 4'b0000;
	mem[3907] = 4'b0000;
	mem[3908] = 4'b0000;
	mem[3909] = 4'b0000;
	mem[3910] = 4'b0001;
	mem[3911] = 4'b1100;
	mem[3912] = 4'b1111;
	mem[3913] = 4'b1111;
	mem[3914] = 4'b1111;
	mem[3915] = 4'b1111;
	mem[3916] = 4'b1101;
	mem[3917] = 4'b1101;
	mem[3918] = 4'b1110;
	mem[3919] = 4'b1111;
	mem[3920] = 4'b1111;
	mem[3921] = 4'b1111;
	mem[3922] = 4'b1111;
	mem[3923] = 4'b1111;
	mem[3924] = 4'b1111;
	mem[3925] = 4'b1111;
	mem[3926] = 4'b1111;
	mem[3927] = 4'b1111;
	mem[3928] = 4'b0100;
	mem[3929] = 4'b0000;
	mem[3930] = 4'b0000;
	mem[3931] = 4'b0000;
	mem[3932] = 4'b0000;
	mem[3933] = 4'b0000;
	mem[3934] = 4'b0000;
	mem[3935] = 4'b0000;
	mem[3936] = 4'b0000;
	mem[3937] = 4'b0000;
	mem[3938] = 4'b0000;
	mem[3939] = 4'b0000;
	mem[3940] = 4'b0000;
	mem[3941] = 4'b0000;
	mem[3942] = 4'b0000;
	mem[3943] = 4'b0000;
	mem[3944] = 4'b0000;
	mem[3945] = 4'b1010;
	mem[3946] = 4'b1111;
	mem[3947] = 4'b1111;
	mem[3948] = 4'b1111;
	mem[3949] = 4'b1111;
	mem[3950] = 4'b1111;
	mem[3951] = 4'b1111;
	mem[3952] = 4'b1111;
	mem[3953] = 4'b1101;
	mem[3954] = 4'b1101;
	mem[3955] = 4'b1110;
	mem[3956] = 4'b1111;
	mem[3957] = 4'b1111;
	mem[3958] = 4'b1111;
	mem[3959] = 4'b1110;
	mem[3960] = 4'b1110;
	mem[3961] = 4'b1110;
	mem[3962] = 4'b0100;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b0111;
	mem[3972] = 4'b1011;
	mem[3973] = 4'b1100;
	mem[3974] = 4'b1110;
	mem[3975] = 4'b1110;
	mem[3976] = 4'b1110;
	mem[3977] = 4'b1101;
	mem[3978] = 4'b1100;
	mem[3979] = 4'b1100;
	mem[3980] = 4'b1110;
	mem[3981] = 4'b1110;
	mem[3982] = 4'b1110;
	mem[3983] = 4'b1110;
	mem[3984] = 4'b1101;
	mem[3985] = 4'b1100;
	mem[3986] = 4'b1100;
	mem[3987] = 4'b1110;
	mem[3988] = 4'b1000;
	mem[3989] = 4'b0110;
	mem[3990] = 4'b0110;
	mem[3991] = 4'b0110;
	mem[3992] = 4'b0110;
	mem[3993] = 4'b0110;
	mem[3994] = 4'b0110;
	mem[3995] = 4'b0011;
	mem[3996] = 4'b0000;
	mem[3997] = 4'b0000;
	mem[3998] = 4'b0000;
	mem[3999] = 4'b0000;
	mem[4000] = 4'b0000;
	mem[4001] = 4'b0000;
	mem[4002] = 4'b0000;
	mem[4003] = 4'b0000;
	mem[4004] = 4'b0000;
	mem[4005] = 4'b1100;
	mem[4006] = 4'b1111;
	mem[4007] = 4'b1111;
	mem[4008] = 4'b1111;
	mem[4009] = 4'b1111;
	mem[4010] = 4'b1111;
	mem[4011] = 4'b1111;
	mem[4012] = 4'b1111;
	mem[4013] = 4'b1111;
	mem[4014] = 4'b1111;
	mem[4015] = 4'b1111;
	mem[4016] = 4'b1111;
	mem[4017] = 4'b1111;
	mem[4018] = 4'b1111;
	mem[4019] = 4'b1111;
	mem[4020] = 4'b1111;
	mem[4021] = 4'b1111;
	mem[4022] = 4'b0110;
	mem[4023] = 4'b0000;
	mem[4024] = 4'b0000;
	mem[4025] = 4'b0000;
	mem[4026] = 4'b0000;
	mem[4027] = 4'b0000;
	mem[4028] = 4'b0000;
	mem[4029] = 4'b0000;
	mem[4030] = 4'b0000;
	mem[4031] = 4'b0000;
	mem[4032] = 4'b0000;
	mem[4033] = 4'b0000;
	mem[4034] = 4'b0000;
	mem[4035] = 4'b0000;
	mem[4036] = 4'b0000;
	mem[4037] = 4'b0001;
	mem[4038] = 4'b0000;
	mem[4039] = 4'b1100;
	mem[4040] = 4'b1111;
	mem[4041] = 4'b1111;
	mem[4042] = 4'b1111;
	mem[4043] = 4'b1111;
	mem[4044] = 4'b1111;
	mem[4045] = 4'b1110;
	mem[4046] = 4'b1111;
	mem[4047] = 4'b1111;
	mem[4048] = 4'b1111;
	mem[4049] = 4'b1111;
	mem[4050] = 4'b1111;
	mem[4051] = 4'b1111;
	mem[4052] = 4'b1111;
	mem[4053] = 4'b1111;
	mem[4054] = 4'b1111;
	mem[4055] = 4'b1111;
	mem[4056] = 4'b0100;
	mem[4057] = 4'b0000;
	mem[4058] = 4'b0000;
	mem[4059] = 4'b0000;
	mem[4060] = 4'b0000;
	mem[4061] = 4'b0000;
	mem[4062] = 4'b0000;
	mem[4063] = 4'b0000;
	mem[4064] = 4'b0000;
	mem[4065] = 4'b0000;
	mem[4066] = 4'b0000;
	mem[4067] = 4'b0000;
	mem[4068] = 4'b0000;
	mem[4069] = 4'b0000;
	mem[4070] = 4'b0000;
	mem[4071] = 4'b0000;
	mem[4072] = 4'b0000;
	mem[4073] = 4'b1010;
	mem[4074] = 4'b1111;
	mem[4075] = 4'b1111;
	mem[4076] = 4'b1111;
	mem[4077] = 4'b1110;
	mem[4078] = 4'b1111;
	mem[4079] = 4'b1111;
	mem[4080] = 4'b1111;
	mem[4081] = 4'b1111;
	mem[4082] = 4'b1101;
	mem[4083] = 4'b1101;
	mem[4084] = 4'b1110;
	mem[4085] = 4'b1110;
	mem[4086] = 4'b1110;
	mem[4087] = 4'b1101;
	mem[4088] = 4'b1111;
	mem[4089] = 4'b1111;
	mem[4090] = 4'b0011;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_2b (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0111;
	mem[4] = 4'b1011;
	mem[5] = 4'b1011;
	mem[6] = 4'b1101;
	mem[7] = 4'b1110;
	mem[8] = 4'b1110;
	mem[9] = 4'b1110;
	mem[10] = 4'b1100;
	mem[11] = 4'b1100;
	mem[12] = 4'b1101;
	mem[13] = 4'b1110;
	mem[14] = 4'b1110;
	mem[15] = 4'b1110;
	mem[16] = 4'b1101;
	mem[17] = 4'b1100;
	mem[18] = 4'b1100;
	mem[19] = 4'b1110;
	mem[20] = 4'b1000;
	mem[21] = 4'b0110;
	mem[22] = 4'b0110;
	mem[23] = 4'b0110;
	mem[24] = 4'b0110;
	mem[25] = 4'b0100;
	mem[26] = 4'b0001;
	mem[27] = 4'b0000;
	mem[28] = 4'b0000;
	mem[29] = 4'b0000;
	mem[30] = 4'b0000;
	mem[31] = 4'b0000;
	mem[32] = 4'b0000;
	mem[33] = 4'b0000;
	mem[34] = 4'b0000;
	mem[35] = 4'b0000;
	mem[36] = 4'b0000;
	mem[37] = 4'b1100;
	mem[38] = 4'b1111;
	mem[39] = 4'b1111;
	mem[40] = 4'b1111;
	mem[41] = 4'b1111;
	mem[42] = 4'b1111;
	mem[43] = 4'b1111;
	mem[44] = 4'b1111;
	mem[45] = 4'b1111;
	mem[46] = 4'b1111;
	mem[47] = 4'b1111;
	mem[48] = 4'b1111;
	mem[49] = 4'b1111;
	mem[50] = 4'b1111;
	mem[51] = 4'b1111;
	mem[52] = 4'b1111;
	mem[53] = 4'b1111;
	mem[54] = 4'b0110;
	mem[55] = 4'b0000;
	mem[56] = 4'b0000;
	mem[57] = 4'b0000;
	mem[58] = 4'b0000;
	mem[59] = 4'b0000;
	mem[60] = 4'b0000;
	mem[61] = 4'b0000;
	mem[62] = 4'b0000;
	mem[63] = 4'b0000;
	mem[64] = 4'b0000;
	mem[65] = 4'b0000;
	mem[66] = 4'b0000;
	mem[67] = 4'b0000;
	mem[68] = 4'b0001;
	mem[69] = 4'b0000;
	mem[70] = 4'b0000;
	mem[71] = 4'b1100;
	mem[72] = 4'b1111;
	mem[73] = 4'b1111;
	mem[74] = 4'b1111;
	mem[75] = 4'b1111;
	mem[76] = 4'b1111;
	mem[77] = 4'b1111;
	mem[78] = 4'b1111;
	mem[79] = 4'b1111;
	mem[80] = 4'b1111;
	mem[81] = 4'b1111;
	mem[82] = 4'b1111;
	mem[83] = 4'b1111;
	mem[84] = 4'b1111;
	mem[85] = 4'b1111;
	mem[86] = 4'b1111;
	mem[87] = 4'b1111;
	mem[88] = 4'b0100;
	mem[89] = 4'b0000;
	mem[90] = 4'b0000;
	mem[91] = 4'b0000;
	mem[92] = 4'b0000;
	mem[93] = 4'b0000;
	mem[94] = 4'b0000;
	mem[95] = 4'b0000;
	mem[96] = 4'b0000;
	mem[97] = 4'b0000;
	mem[98] = 4'b0000;
	mem[99] = 4'b0000;
	mem[100] = 4'b0000;
	mem[101] = 4'b0000;
	mem[102] = 4'b0000;
	mem[103] = 4'b0000;
	mem[104] = 4'b0000;
	mem[105] = 4'b1010;
	mem[106] = 4'b1111;
	mem[107] = 4'b1110;
	mem[108] = 4'b1101;
	mem[109] = 4'b1101;
	mem[110] = 4'b1101;
	mem[111] = 4'b1110;
	mem[112] = 4'b1111;
	mem[113] = 4'b1111;
	mem[114] = 4'b1111;
	mem[115] = 4'b1101;
	mem[116] = 4'b1101;
	mem[117] = 4'b1101;
	mem[118] = 4'b1101;
	mem[119] = 4'b1110;
	mem[120] = 4'b1111;
	mem[121] = 4'b1111;
	mem[122] = 4'b0011;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b1000;
	mem[132] = 4'b1100;
	mem[133] = 4'b1011;
	mem[134] = 4'b1100;
	mem[135] = 4'b1101;
	mem[136] = 4'b1110;
	mem[137] = 4'b1110;
	mem[138] = 4'b1101;
	mem[139] = 4'b1100;
	mem[140] = 4'b1100;
	mem[141] = 4'b1101;
	mem[142] = 4'b1101;
	mem[143] = 4'b1101;
	mem[144] = 4'b1100;
	mem[145] = 4'b1100;
	mem[146] = 4'b1101;
	mem[147] = 4'b1110;
	mem[148] = 4'b1000;
	mem[149] = 4'b0110;
	mem[150] = 4'b0110;
	mem[151] = 4'b0110;
	mem[152] = 4'b0010;
	mem[153] = 4'b0000;
	mem[154] = 4'b0000;
	mem[155] = 4'b0000;
	mem[156] = 4'b0000;
	mem[157] = 4'b0000;
	mem[158] = 4'b0000;
	mem[159] = 4'b0000;
	mem[160] = 4'b0000;
	mem[161] = 4'b0000;
	mem[162] = 4'b0000;
	mem[163] = 4'b0000;
	mem[164] = 4'b0000;
	mem[165] = 4'b1100;
	mem[166] = 4'b1111;
	mem[167] = 4'b1111;
	mem[168] = 4'b1111;
	mem[169] = 4'b1111;
	mem[170] = 4'b1111;
	mem[171] = 4'b1111;
	mem[172] = 4'b1111;
	mem[173] = 4'b1111;
	mem[174] = 4'b1111;
	mem[175] = 4'b1111;
	mem[176] = 4'b1111;
	mem[177] = 4'b1111;
	mem[178] = 4'b1111;
	mem[179] = 4'b1111;
	mem[180] = 4'b1111;
	mem[181] = 4'b1111;
	mem[182] = 4'b0101;
	mem[183] = 4'b0000;
	mem[184] = 4'b0000;
	mem[185] = 4'b0000;
	mem[186] = 4'b0000;
	mem[187] = 4'b0000;
	mem[188] = 4'b0000;
	mem[189] = 4'b0000;
	mem[190] = 4'b0000;
	mem[191] = 4'b0000;
	mem[192] = 4'b0000;
	mem[193] = 4'b0000;
	mem[194] = 4'b0000;
	mem[195] = 4'b0001;
	mem[196] = 4'b0000;
	mem[197] = 4'b0000;
	mem[198] = 4'b0000;
	mem[199] = 4'b1100;
	mem[200] = 4'b1111;
	mem[201] = 4'b1111;
	mem[202] = 4'b1111;
	mem[203] = 4'b1111;
	mem[204] = 4'b1111;
	mem[205] = 4'b1111;
	mem[206] = 4'b1111;
	mem[207] = 4'b1111;
	mem[208] = 4'b1111;
	mem[209] = 4'b1111;
	mem[210] = 4'b1111;
	mem[211] = 4'b1111;
	mem[212] = 4'b1111;
	mem[213] = 4'b1111;
	mem[214] = 4'b1111;
	mem[215] = 4'b1111;
	mem[216] = 4'b0100;
	mem[217] = 4'b0000;
	mem[218] = 4'b0000;
	mem[219] = 4'b0000;
	mem[220] = 4'b0000;
	mem[221] = 4'b0000;
	mem[222] = 4'b0000;
	mem[223] = 4'b0000;
	mem[224] = 4'b0000;
	mem[225] = 4'b0000;
	mem[226] = 4'b0000;
	mem[227] = 4'b0000;
	mem[228] = 4'b0000;
	mem[229] = 4'b0000;
	mem[230] = 4'b0000;
	mem[231] = 4'b0000;
	mem[232] = 4'b0000;
	mem[233] = 4'b1010;
	mem[234] = 4'b1111;
	mem[235] = 4'b1101;
	mem[236] = 4'b1110;
	mem[237] = 4'b1110;
	mem[238] = 4'b1101;
	mem[239] = 4'b1101;
	mem[240] = 4'b1110;
	mem[241] = 4'b1111;
	mem[242] = 4'b1111;
	mem[243] = 4'b1111;
	mem[244] = 4'b1111;
	mem[245] = 4'b1111;
	mem[246] = 4'b1111;
	mem[247] = 4'b1111;
	mem[248] = 4'b1111;
	mem[249] = 4'b1111;
	mem[250] = 4'b0011;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0111;
	mem[260] = 4'b1100;
	mem[261] = 4'b1100;
	mem[262] = 4'b1100;
	mem[263] = 4'b1100;
	mem[264] = 4'b1101;
	mem[265] = 4'b1110;
	mem[266] = 4'b1110;
	mem[267] = 4'b1101;
	mem[268] = 4'b1100;
	mem[269] = 4'b1100;
	mem[270] = 4'b1100;
	mem[271] = 4'b1100;
	mem[272] = 4'b1100;
	mem[273] = 4'b1101;
	mem[274] = 4'b1110;
	mem[275] = 4'b1110;
	mem[276] = 4'b1000;
	mem[277] = 4'b0110;
	mem[278] = 4'b0011;
	mem[279] = 4'b0000;
	mem[280] = 4'b0000;
	mem[281] = 4'b0000;
	mem[282] = 4'b0000;
	mem[283] = 4'b0000;
	mem[284] = 4'b0000;
	mem[285] = 4'b0000;
	mem[286] = 4'b0000;
	mem[287] = 4'b0000;
	mem[288] = 4'b0000;
	mem[289] = 4'b0000;
	mem[290] = 4'b0000;
	mem[291] = 4'b0000;
	mem[292] = 4'b0000;
	mem[293] = 4'b1100;
	mem[294] = 4'b1111;
	mem[295] = 4'b1111;
	mem[296] = 4'b1111;
	mem[297] = 4'b1111;
	mem[298] = 4'b1111;
	mem[299] = 4'b1111;
	mem[300] = 4'b1111;
	mem[301] = 4'b1111;
	mem[302] = 4'b1111;
	mem[303] = 4'b1111;
	mem[304] = 4'b1111;
	mem[305] = 4'b1111;
	mem[306] = 4'b1111;
	mem[307] = 4'b1111;
	mem[308] = 4'b1110;
	mem[309] = 4'b1101;
	mem[310] = 4'b0101;
	mem[311] = 4'b0000;
	mem[312] = 4'b0000;
	mem[313] = 4'b0000;
	mem[314] = 4'b0001;
	mem[315] = 4'b0000;
	mem[316] = 4'b0000;
	mem[317] = 4'b0000;
	mem[318] = 4'b0000;
	mem[319] = 4'b0000;
	mem[320] = 4'b0000;
	mem[321] = 4'b0000;
	mem[322] = 4'b0001;
	mem[323] = 4'b0000;
	mem[324] = 4'b0000;
	mem[325] = 4'b0000;
	mem[326] = 4'b0000;
	mem[327] = 4'b1100;
	mem[328] = 4'b1111;
	mem[329] = 4'b1111;
	mem[330] = 4'b1111;
	mem[331] = 4'b1111;
	mem[332] = 4'b1111;
	mem[333] = 4'b1111;
	mem[334] = 4'b1111;
	mem[335] = 4'b1111;
	mem[336] = 4'b1111;
	mem[337] = 4'b1111;
	mem[338] = 4'b1111;
	mem[339] = 4'b1111;
	mem[340] = 4'b1111;
	mem[341] = 4'b1111;
	mem[342] = 4'b1111;
	mem[343] = 4'b1111;
	mem[344] = 4'b0100;
	mem[345] = 4'b0000;
	mem[346] = 4'b0000;
	mem[347] = 4'b0000;
	mem[348] = 4'b0000;
	mem[349] = 4'b0000;
	mem[350] = 4'b0000;
	mem[351] = 4'b0000;
	mem[352] = 4'b0000;
	mem[353] = 4'b0000;
	mem[354] = 4'b0000;
	mem[355] = 4'b0000;
	mem[356] = 4'b0000;
	mem[357] = 4'b0000;
	mem[358] = 4'b0000;
	mem[359] = 4'b0000;
	mem[360] = 4'b0000;
	mem[361] = 4'b1001;
	mem[362] = 4'b1110;
	mem[363] = 4'b1110;
	mem[364] = 4'b1111;
	mem[365] = 4'b1111;
	mem[366] = 4'b1111;
	mem[367] = 4'b1101;
	mem[368] = 4'b1101;
	mem[369] = 4'b1110;
	mem[370] = 4'b1111;
	mem[371] = 4'b1111;
	mem[372] = 4'b1111;
	mem[373] = 4'b1111;
	mem[374] = 4'b1111;
	mem[375] = 4'b1111;
	mem[376] = 4'b1111;
	mem[377] = 4'b1111;
	mem[378] = 4'b0011;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0111;
	mem[388] = 4'b1100;
	mem[389] = 4'b1101;
	mem[390] = 4'b1101;
	mem[391] = 4'b1100;
	mem[392] = 4'b1100;
	mem[393] = 4'b1101;
	mem[394] = 4'b1110;
	mem[395] = 4'b1110;
	mem[396] = 4'b1101;
	mem[397] = 4'b1100;
	mem[398] = 4'b1100;
	mem[399] = 4'b1100;
	mem[400] = 4'b1101;
	mem[401] = 4'b1110;
	mem[402] = 4'b1110;
	mem[403] = 4'b1110;
	mem[404] = 4'b0111;
	mem[405] = 4'b0001;
	mem[406] = 4'b0000;
	mem[407] = 4'b0000;
	mem[408] = 4'b0000;
	mem[409] = 4'b0000;
	mem[410] = 4'b0000;
	mem[411] = 4'b0000;
	mem[412] = 4'b0000;
	mem[413] = 4'b0000;
	mem[414] = 4'b0000;
	mem[415] = 4'b0000;
	mem[416] = 4'b0000;
	mem[417] = 4'b0000;
	mem[418] = 4'b0000;
	mem[419] = 4'b0000;
	mem[420] = 4'b0000;
	mem[421] = 4'b1100;
	mem[422] = 4'b1111;
	mem[423] = 4'b1111;
	mem[424] = 4'b1111;
	mem[425] = 4'b1111;
	mem[426] = 4'b1111;
	mem[427] = 4'b1111;
	mem[428] = 4'b1111;
	mem[429] = 4'b1111;
	mem[430] = 4'b1111;
	mem[431] = 4'b1111;
	mem[432] = 4'b1111;
	mem[433] = 4'b1111;
	mem[434] = 4'b1111;
	mem[435] = 4'b1110;
	mem[436] = 4'b1101;
	mem[437] = 4'b1101;
	mem[438] = 4'b0101;
	mem[439] = 4'b0000;
	mem[440] = 4'b0000;
	mem[441] = 4'b0001;
	mem[442] = 4'b0001;
	mem[443] = 4'b0000;
	mem[444] = 4'b0000;
	mem[445] = 4'b0000;
	mem[446] = 4'b0000;
	mem[447] = 4'b0000;
	mem[448] = 4'b0000;
	mem[449] = 4'b0000;
	mem[450] = 4'b0000;
	mem[451] = 4'b0000;
	mem[452] = 4'b0000;
	mem[453] = 4'b0000;
	mem[454] = 4'b0000;
	mem[455] = 4'b1100;
	mem[456] = 4'b1111;
	mem[457] = 4'b1111;
	mem[458] = 4'b1111;
	mem[459] = 4'b1111;
	mem[460] = 4'b1111;
	mem[461] = 4'b1111;
	mem[462] = 4'b1111;
	mem[463] = 4'b1111;
	mem[464] = 4'b1111;
	mem[465] = 4'b1111;
	mem[466] = 4'b1111;
	mem[467] = 4'b1111;
	mem[468] = 4'b1111;
	mem[469] = 4'b1111;
	mem[470] = 4'b1111;
	mem[471] = 4'b1111;
	mem[472] = 4'b0100;
	mem[473] = 4'b0000;
	mem[474] = 4'b0000;
	mem[475] = 4'b0000;
	mem[476] = 4'b0000;
	mem[477] = 4'b0000;
	mem[478] = 4'b0000;
	mem[479] = 4'b0000;
	mem[480] = 4'b0000;
	mem[481] = 4'b0000;
	mem[482] = 4'b0000;
	mem[483] = 4'b0000;
	mem[484] = 4'b0000;
	mem[485] = 4'b0000;
	mem[486] = 4'b0000;
	mem[487] = 4'b0000;
	mem[488] = 4'b0000;
	mem[489] = 4'b1000;
	mem[490] = 4'b1101;
	mem[491] = 4'b1111;
	mem[492] = 4'b1111;
	mem[493] = 4'b1111;
	mem[494] = 4'b1111;
	mem[495] = 4'b1111;
	mem[496] = 4'b1101;
	mem[497] = 4'b1101;
	mem[498] = 4'b1110;
	mem[499] = 4'b1111;
	mem[500] = 4'b1111;
	mem[501] = 4'b1111;
	mem[502] = 4'b1111;
	mem[503] = 4'b1111;
	mem[504] = 4'b1111;
	mem[505] = 4'b1111;
	mem[506] = 4'b0011;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0111;
	mem[516] = 4'b1100;
	mem[517] = 4'b1101;
	mem[518] = 4'b1110;
	mem[519] = 4'b1101;
	mem[520] = 4'b1100;
	mem[521] = 4'b1100;
	mem[522] = 4'b1101;
	mem[523] = 4'b1110;
	mem[524] = 4'b1110;
	mem[525] = 4'b1110;
	mem[526] = 4'b1110;
	mem[527] = 4'b1110;
	mem[528] = 4'b1110;
	mem[529] = 4'b1110;
	mem[530] = 4'b1110;
	mem[531] = 4'b1101;
	mem[532] = 4'b0011;
	mem[533] = 4'b0000;
	mem[534] = 4'b0000;
	mem[535] = 4'b0000;
	mem[536] = 4'b0000;
	mem[537] = 4'b0000;
	mem[538] = 4'b0000;
	mem[539] = 4'b0000;
	mem[540] = 4'b0000;
	mem[541] = 4'b0000;
	mem[542] = 4'b0000;
	mem[543] = 4'b0000;
	mem[544] = 4'b0000;
	mem[545] = 4'b0000;
	mem[546] = 4'b0000;
	mem[547] = 4'b0000;
	mem[548] = 4'b0000;
	mem[549] = 4'b1100;
	mem[550] = 4'b1111;
	mem[551] = 4'b1111;
	mem[552] = 4'b1111;
	mem[553] = 4'b1111;
	mem[554] = 4'b1111;
	mem[555] = 4'b1111;
	mem[556] = 4'b1111;
	mem[557] = 4'b1111;
	mem[558] = 4'b1111;
	mem[559] = 4'b1111;
	mem[560] = 4'b1111;
	mem[561] = 4'b1111;
	mem[562] = 4'b1110;
	mem[563] = 4'b1101;
	mem[564] = 4'b1101;
	mem[565] = 4'b1101;
	mem[566] = 4'b0110;
	mem[567] = 4'b0001;
	mem[568] = 4'b0001;
	mem[569] = 4'b0001;
	mem[570] = 4'b0000;
	mem[571] = 4'b0000;
	mem[572] = 4'b0000;
	mem[573] = 4'b0000;
	mem[574] = 4'b0000;
	mem[575] = 4'b0000;
	mem[576] = 4'b0000;
	mem[577] = 4'b0000;
	mem[578] = 4'b0000;
	mem[579] = 4'b0000;
	mem[580] = 4'b0000;
	mem[581] = 4'b0000;
	mem[582] = 4'b0000;
	mem[583] = 4'b1100;
	mem[584] = 4'b1111;
	mem[585] = 4'b1111;
	mem[586] = 4'b1111;
	mem[587] = 4'b1111;
	mem[588] = 4'b1111;
	mem[589] = 4'b1111;
	mem[590] = 4'b1111;
	mem[591] = 4'b1111;
	mem[592] = 4'b1111;
	mem[593] = 4'b1111;
	mem[594] = 4'b1111;
	mem[595] = 4'b1111;
	mem[596] = 4'b1111;
	mem[597] = 4'b1111;
	mem[598] = 4'b1111;
	mem[599] = 4'b1111;
	mem[600] = 4'b0100;
	mem[601] = 4'b0000;
	mem[602] = 4'b0000;
	mem[603] = 4'b0000;
	mem[604] = 4'b0000;
	mem[605] = 4'b0000;
	mem[606] = 4'b0000;
	mem[607] = 4'b0000;
	mem[608] = 4'b0000;
	mem[609] = 4'b0000;
	mem[610] = 4'b0000;
	mem[611] = 4'b0000;
	mem[612] = 4'b0000;
	mem[613] = 4'b0000;
	mem[614] = 4'b0000;
	mem[615] = 4'b0000;
	mem[616] = 4'b0000;
	mem[617] = 4'b1000;
	mem[618] = 4'b1101;
	mem[619] = 4'b1110;
	mem[620] = 4'b1111;
	mem[621] = 4'b1111;
	mem[622] = 4'b1111;
	mem[623] = 4'b1111;
	mem[624] = 4'b1111;
	mem[625] = 4'b1101;
	mem[626] = 4'b1101;
	mem[627] = 4'b1111;
	mem[628] = 4'b1111;
	mem[629] = 4'b1111;
	mem[630] = 4'b1111;
	mem[631] = 4'b1111;
	mem[632] = 4'b1111;
	mem[633] = 4'b1111;
	mem[634] = 4'b0011;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0111;
	mem[644] = 4'b1100;
	mem[645] = 4'b1101;
	mem[646] = 4'b1110;
	mem[647] = 4'b1110;
	mem[648] = 4'b1101;
	mem[649] = 4'b1100;
	mem[650] = 4'b1100;
	mem[651] = 4'b1101;
	mem[652] = 4'b1110;
	mem[653] = 4'b1110;
	mem[654] = 4'b1110;
	mem[655] = 4'b1110;
	mem[656] = 4'b1110;
	mem[657] = 4'b1101;
	mem[658] = 4'b1100;
	mem[659] = 4'b1100;
	mem[660] = 4'b0011;
	mem[661] = 4'b0000;
	mem[662] = 4'b0000;
	mem[663] = 4'b0000;
	mem[664] = 4'b0000;
	mem[665] = 4'b0000;
	mem[666] = 4'b0000;
	mem[667] = 4'b0000;
	mem[668] = 4'b0000;
	mem[669] = 4'b0000;
	mem[670] = 4'b0000;
	mem[671] = 4'b0000;
	mem[672] = 4'b0000;
	mem[673] = 4'b0000;
	mem[674] = 4'b0000;
	mem[675] = 4'b0000;
	mem[676] = 4'b0000;
	mem[677] = 4'b1100;
	mem[678] = 4'b1111;
	mem[679] = 4'b1111;
	mem[680] = 4'b1111;
	mem[681] = 4'b1111;
	mem[682] = 4'b1111;
	mem[683] = 4'b1111;
	mem[684] = 4'b1111;
	mem[685] = 4'b1111;
	mem[686] = 4'b1111;
	mem[687] = 4'b1111;
	mem[688] = 4'b1111;
	mem[689] = 4'b1111;
	mem[690] = 4'b1101;
	mem[691] = 4'b1101;
	mem[692] = 4'b1101;
	mem[693] = 4'b1111;
	mem[694] = 4'b0110;
	mem[695] = 4'b0000;
	mem[696] = 4'b0000;
	mem[697] = 4'b0000;
	mem[698] = 4'b0000;
	mem[699] = 4'b0000;
	mem[700] = 4'b0000;
	mem[701] = 4'b0000;
	mem[702] = 4'b0000;
	mem[703] = 4'b0000;
	mem[704] = 4'b0000;
	mem[705] = 4'b0000;
	mem[706] = 4'b0000;
	mem[707] = 4'b0000;
	mem[708] = 4'b0000;
	mem[709] = 4'b0000;
	mem[710] = 4'b0000;
	mem[711] = 4'b1100;
	mem[712] = 4'b1111;
	mem[713] = 4'b1111;
	mem[714] = 4'b1111;
	mem[715] = 4'b1111;
	mem[716] = 4'b1111;
	mem[717] = 4'b1111;
	mem[718] = 4'b1111;
	mem[719] = 4'b1111;
	mem[720] = 4'b1111;
	mem[721] = 4'b1111;
	mem[722] = 4'b1111;
	mem[723] = 4'b1111;
	mem[724] = 4'b1111;
	mem[725] = 4'b1111;
	mem[726] = 4'b1111;
	mem[727] = 4'b1111;
	mem[728] = 4'b0100;
	mem[729] = 4'b0000;
	mem[730] = 4'b0000;
	mem[731] = 4'b0000;
	mem[732] = 4'b0000;
	mem[733] = 4'b0000;
	mem[734] = 4'b0000;
	mem[735] = 4'b0000;
	mem[736] = 4'b0000;
	mem[737] = 4'b0000;
	mem[738] = 4'b0000;
	mem[739] = 4'b0000;
	mem[740] = 4'b0000;
	mem[741] = 4'b0000;
	mem[742] = 4'b0000;
	mem[743] = 4'b0000;
	mem[744] = 4'b0000;
	mem[745] = 4'b1001;
	mem[746] = 4'b1101;
	mem[747] = 4'b1101;
	mem[748] = 4'b1110;
	mem[749] = 4'b1111;
	mem[750] = 4'b1111;
	mem[751] = 4'b1111;
	mem[752] = 4'b1111;
	mem[753] = 4'b1111;
	mem[754] = 4'b1110;
	mem[755] = 4'b1111;
	mem[756] = 4'b1111;
	mem[757] = 4'b1111;
	mem[758] = 4'b1111;
	mem[759] = 4'b1111;
	mem[760] = 4'b1111;
	mem[761] = 4'b1111;
	mem[762] = 4'b0011;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0111;
	mem[772] = 4'b1100;
	mem[773] = 4'b1101;
	mem[774] = 4'b1110;
	mem[775] = 4'b1110;
	mem[776] = 4'b1110;
	mem[777] = 4'b1101;
	mem[778] = 4'b1100;
	mem[779] = 4'b1100;
	mem[780] = 4'b1101;
	mem[781] = 4'b1110;
	mem[782] = 4'b1110;
	mem[783] = 4'b1110;
	mem[784] = 4'b1101;
	mem[785] = 4'b1100;
	mem[786] = 4'b1100;
	mem[787] = 4'b1100;
	mem[788] = 4'b0011;
	mem[789] = 4'b0000;
	mem[790] = 4'b0000;
	mem[791] = 4'b0000;
	mem[792] = 4'b0000;
	mem[793] = 4'b0000;
	mem[794] = 4'b0000;
	mem[795] = 4'b0000;
	mem[796] = 4'b0000;
	mem[797] = 4'b0000;
	mem[798] = 4'b0000;
	mem[799] = 4'b0000;
	mem[800] = 4'b0000;
	mem[801] = 4'b0000;
	mem[802] = 4'b0000;
	mem[803] = 4'b0000;
	mem[804] = 4'b0000;
	mem[805] = 4'b1100;
	mem[806] = 4'b1111;
	mem[807] = 4'b1111;
	mem[808] = 4'b1111;
	mem[809] = 4'b1111;
	mem[810] = 4'b1111;
	mem[811] = 4'b1111;
	mem[812] = 4'b1111;
	mem[813] = 4'b1111;
	mem[814] = 4'b1111;
	mem[815] = 4'b1111;
	mem[816] = 4'b1111;
	mem[817] = 4'b1110;
	mem[818] = 4'b1101;
	mem[819] = 4'b1101;
	mem[820] = 4'b1110;
	mem[821] = 4'b1111;
	mem[822] = 4'b0110;
	mem[823] = 4'b0000;
	mem[824] = 4'b0000;
	mem[825] = 4'b0000;
	mem[826] = 4'b0000;
	mem[827] = 4'b0000;
	mem[828] = 4'b0000;
	mem[829] = 4'b0000;
	mem[830] = 4'b0000;
	mem[831] = 4'b0000;
	mem[832] = 4'b0000;
	mem[833] = 4'b0000;
	mem[834] = 4'b0000;
	mem[835] = 4'b0000;
	mem[836] = 4'b0000;
	mem[837] = 4'b0000;
	mem[838] = 4'b0000;
	mem[839] = 4'b1100;
	mem[840] = 4'b1111;
	mem[841] = 4'b1111;
	mem[842] = 4'b1111;
	mem[843] = 4'b1111;
	mem[844] = 4'b1111;
	mem[845] = 4'b1111;
	mem[846] = 4'b1111;
	mem[847] = 4'b1111;
	mem[848] = 4'b1111;
	mem[849] = 4'b1111;
	mem[850] = 4'b1111;
	mem[851] = 4'b1111;
	mem[852] = 4'b1111;
	mem[853] = 4'b1111;
	mem[854] = 4'b1111;
	mem[855] = 4'b1111;
	mem[856] = 4'b0100;
	mem[857] = 4'b0000;
	mem[858] = 4'b0000;
	mem[859] = 4'b0000;
	mem[860] = 4'b0000;
	mem[861] = 4'b0000;
	mem[862] = 4'b0000;
	mem[863] = 4'b0000;
	mem[864] = 4'b0000;
	mem[865] = 4'b0000;
	mem[866] = 4'b0000;
	mem[867] = 4'b0000;
	mem[868] = 4'b0000;
	mem[869] = 4'b0000;
	mem[870] = 4'b0000;
	mem[871] = 4'b0000;
	mem[872] = 4'b0000;
	mem[873] = 4'b1010;
	mem[874] = 4'b1111;
	mem[875] = 4'b1101;
	mem[876] = 4'b1101;
	mem[877] = 4'b1110;
	mem[878] = 4'b1111;
	mem[879] = 4'b1111;
	mem[880] = 4'b1111;
	mem[881] = 4'b1111;
	mem[882] = 4'b1111;
	mem[883] = 4'b1111;
	mem[884] = 4'b1111;
	mem[885] = 4'b1111;
	mem[886] = 4'b1111;
	mem[887] = 4'b1111;
	mem[888] = 4'b1111;
	mem[889] = 4'b1111;
	mem[890] = 4'b0011;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0111;
	mem[900] = 4'b1100;
	mem[901] = 4'b1101;
	mem[902] = 4'b1110;
	mem[903] = 4'b1110;
	mem[904] = 4'b1110;
	mem[905] = 4'b1110;
	mem[906] = 4'b1101;
	mem[907] = 4'b1100;
	mem[908] = 4'b1101;
	mem[909] = 4'b1110;
	mem[910] = 4'b1101;
	mem[911] = 4'b1101;
	mem[912] = 4'b1100;
	mem[913] = 4'b1100;
	mem[914] = 4'b1100;
	mem[915] = 4'b1100;
	mem[916] = 4'b0011;
	mem[917] = 4'b0000;
	mem[918] = 4'b0000;
	mem[919] = 4'b0000;
	mem[920] = 4'b0000;
	mem[921] = 4'b0000;
	mem[922] = 4'b0000;
	mem[923] = 4'b0000;
	mem[924] = 4'b0000;
	mem[925] = 4'b0000;
	mem[926] = 4'b0000;
	mem[927] = 4'b0000;
	mem[928] = 4'b0000;
	mem[929] = 4'b0000;
	mem[930] = 4'b0000;
	mem[931] = 4'b0000;
	mem[932] = 4'b0000;
	mem[933] = 4'b1100;
	mem[934] = 4'b1111;
	mem[935] = 4'b1111;
	mem[936] = 4'b1111;
	mem[937] = 4'b1111;
	mem[938] = 4'b1111;
	mem[939] = 4'b1111;
	mem[940] = 4'b1111;
	mem[941] = 4'b1111;
	mem[942] = 4'b1111;
	mem[943] = 4'b1111;
	mem[944] = 4'b1111;
	mem[945] = 4'b1110;
	mem[946] = 4'b1101;
	mem[947] = 4'b1101;
	mem[948] = 4'b1111;
	mem[949] = 4'b1111;
	mem[950] = 4'b0101;
	mem[951] = 4'b0000;
	mem[952] = 4'b0000;
	mem[953] = 4'b0000;
	mem[954] = 4'b0000;
	mem[955] = 4'b0000;
	mem[956] = 4'b0000;
	mem[957] = 4'b0000;
	mem[958] = 4'b0000;
	mem[959] = 4'b0000;
	mem[960] = 4'b0000;
	mem[961] = 4'b0001;
	mem[962] = 4'b0000;
	mem[963] = 4'b0000;
	mem[964] = 4'b0000;
	mem[965] = 4'b0000;
	mem[966] = 4'b0000;
	mem[967] = 4'b1100;
	mem[968] = 4'b1111;
	mem[969] = 4'b1111;
	mem[970] = 4'b1111;
	mem[971] = 4'b1111;
	mem[972] = 4'b1111;
	mem[973] = 4'b1111;
	mem[974] = 4'b1111;
	mem[975] = 4'b1111;
	mem[976] = 4'b1111;
	mem[977] = 4'b1111;
	mem[978] = 4'b1111;
	mem[979] = 4'b1111;
	mem[980] = 4'b1111;
	mem[981] = 4'b1111;
	mem[982] = 4'b1111;
	mem[983] = 4'b1111;
	mem[984] = 4'b0100;
	mem[985] = 4'b0000;
	mem[986] = 4'b0000;
	mem[987] = 4'b0000;
	mem[988] = 4'b0000;
	mem[989] = 4'b0000;
	mem[990] = 4'b0000;
	mem[991] = 4'b0000;
	mem[992] = 4'b0000;
	mem[993] = 4'b0000;
	mem[994] = 4'b0000;
	mem[995] = 4'b0000;
	mem[996] = 4'b0000;
	mem[997] = 4'b0000;
	mem[998] = 4'b0000;
	mem[999] = 4'b0000;
	mem[1000] = 4'b0000;
	mem[1001] = 4'b1010;
	mem[1002] = 4'b1111;
	mem[1003] = 4'b1111;
	mem[1004] = 4'b1101;
	mem[1005] = 4'b1101;
	mem[1006] = 4'b1110;
	mem[1007] = 4'b1111;
	mem[1008] = 4'b1111;
	mem[1009] = 4'b1111;
	mem[1010] = 4'b1111;
	mem[1011] = 4'b1111;
	mem[1012] = 4'b1111;
	mem[1013] = 4'b1111;
	mem[1014] = 4'b1111;
	mem[1015] = 4'b1111;
	mem[1016] = 4'b1111;
	mem[1017] = 4'b1111;
	mem[1018] = 4'b0011;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0111;
	mem[1028] = 4'b1100;
	mem[1029] = 4'b1101;
	mem[1030] = 4'b1110;
	mem[1031] = 4'b1110;
	mem[1032] = 4'b1110;
	mem[1033] = 4'b1110;
	mem[1034] = 4'b1110;
	mem[1035] = 4'b1101;
	mem[1036] = 4'b1110;
	mem[1037] = 4'b1101;
	mem[1038] = 4'b1100;
	mem[1039] = 4'b1100;
	mem[1040] = 4'b1100;
	mem[1041] = 4'b1100;
	mem[1042] = 4'b1100;
	mem[1043] = 4'b1100;
	mem[1044] = 4'b0011;
	mem[1045] = 4'b0000;
	mem[1046] = 4'b0000;
	mem[1047] = 4'b0000;
	mem[1048] = 4'b0000;
	mem[1049] = 4'b0000;
	mem[1050] = 4'b0000;
	mem[1051] = 4'b0000;
	mem[1052] = 4'b0000;
	mem[1053] = 4'b0000;
	mem[1054] = 4'b0000;
	mem[1055] = 4'b0000;
	mem[1056] = 4'b0000;
	mem[1057] = 4'b0000;
	mem[1058] = 4'b0000;
	mem[1059] = 4'b0000;
	mem[1060] = 4'b0000;
	mem[1061] = 4'b1100;
	mem[1062] = 4'b1111;
	mem[1063] = 4'b1111;
	mem[1064] = 4'b1111;
	mem[1065] = 4'b1111;
	mem[1066] = 4'b1111;
	mem[1067] = 4'b1111;
	mem[1068] = 4'b1111;
	mem[1069] = 4'b1111;
	mem[1070] = 4'b1111;
	mem[1071] = 4'b1111;
	mem[1072] = 4'b1111;
	mem[1073] = 4'b1110;
	mem[1074] = 4'b1101;
	mem[1075] = 4'b1101;
	mem[1076] = 4'b1110;
	mem[1077] = 4'b1110;
	mem[1078] = 4'b0101;
	mem[1079] = 4'b0000;
	mem[1080] = 4'b0000;
	mem[1081] = 4'b0000;
	mem[1082] = 4'b0000;
	mem[1083] = 4'b0000;
	mem[1084] = 4'b0001;
	mem[1085] = 4'b0000;
	mem[1086] = 4'b0000;
	mem[1087] = 4'b0000;
	mem[1088] = 4'b0000;
	mem[1089] = 4'b0001;
	mem[1090] = 4'b0000;
	mem[1091] = 4'b0000;
	mem[1092] = 4'b0000;
	mem[1093] = 4'b0000;
	mem[1094] = 4'b0000;
	mem[1095] = 4'b1100;
	mem[1096] = 4'b1111;
	mem[1097] = 4'b1111;
	mem[1098] = 4'b1111;
	mem[1099] = 4'b1111;
	mem[1100] = 4'b1111;
	mem[1101] = 4'b1111;
	mem[1102] = 4'b1111;
	mem[1103] = 4'b1111;
	mem[1104] = 4'b1111;
	mem[1105] = 4'b1111;
	mem[1106] = 4'b1111;
	mem[1107] = 4'b1111;
	mem[1108] = 4'b1111;
	mem[1109] = 4'b1111;
	mem[1110] = 4'b1111;
	mem[1111] = 4'b1111;
	mem[1112] = 4'b0100;
	mem[1113] = 4'b0000;
	mem[1114] = 4'b0000;
	mem[1115] = 4'b0000;
	mem[1116] = 4'b0000;
	mem[1117] = 4'b0000;
	mem[1118] = 4'b0000;
	mem[1119] = 4'b0000;
	mem[1120] = 4'b0000;
	mem[1121] = 4'b0000;
	mem[1122] = 4'b0000;
	mem[1123] = 4'b0000;
	mem[1124] = 4'b0000;
	mem[1125] = 4'b0001;
	mem[1126] = 4'b0000;
	mem[1127] = 4'b0000;
	mem[1128] = 4'b0000;
	mem[1129] = 4'b1001;
	mem[1130] = 4'b1111;
	mem[1131] = 4'b1111;
	mem[1132] = 4'b1111;
	mem[1133] = 4'b1101;
	mem[1134] = 4'b1101;
	mem[1135] = 4'b1111;
	mem[1136] = 4'b1111;
	mem[1137] = 4'b1111;
	mem[1138] = 4'b1111;
	mem[1139] = 4'b1111;
	mem[1140] = 4'b1111;
	mem[1141] = 4'b1111;
	mem[1142] = 4'b1111;
	mem[1143] = 4'b1111;
	mem[1144] = 4'b1111;
	mem[1145] = 4'b1111;
	mem[1146] = 4'b0011;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0111;
	mem[1156] = 4'b1100;
	mem[1157] = 4'b1101;
	mem[1158] = 4'b1110;
	mem[1159] = 4'b1110;
	mem[1160] = 4'b1110;
	mem[1161] = 4'b1110;
	mem[1162] = 4'b1110;
	mem[1163] = 4'b1110;
	mem[1164] = 4'b1101;
	mem[1165] = 4'b1100;
	mem[1166] = 4'b1100;
	mem[1167] = 4'b1100;
	mem[1168] = 4'b1100;
	mem[1169] = 4'b1100;
	mem[1170] = 4'b1100;
	mem[1171] = 4'b1100;
	mem[1172] = 4'b0011;
	mem[1173] = 4'b0000;
	mem[1174] = 4'b0000;
	mem[1175] = 4'b0000;
	mem[1176] = 4'b0000;
	mem[1177] = 4'b0000;
	mem[1178] = 4'b0000;
	mem[1179] = 4'b0000;
	mem[1180] = 4'b0000;
	mem[1181] = 4'b0000;
	mem[1182] = 4'b0000;
	mem[1183] = 4'b0000;
	mem[1184] = 4'b0000;
	mem[1185] = 4'b0000;
	mem[1186] = 4'b0000;
	mem[1187] = 4'b0000;
	mem[1188] = 4'b0000;
	mem[1189] = 4'b1100;
	mem[1190] = 4'b1111;
	mem[1191] = 4'b1111;
	mem[1192] = 4'b1111;
	mem[1193] = 4'b1111;
	mem[1194] = 4'b1111;
	mem[1195] = 4'b1111;
	mem[1196] = 4'b1111;
	mem[1197] = 4'b1111;
	mem[1198] = 4'b1111;
	mem[1199] = 4'b1111;
	mem[1200] = 4'b1111;
	mem[1201] = 4'b1110;
	mem[1202] = 4'b1101;
	mem[1203] = 4'b1101;
	mem[1204] = 4'b1101;
	mem[1205] = 4'b1101;
	mem[1206] = 4'b0101;
	mem[1207] = 4'b0000;
	mem[1208] = 4'b0000;
	mem[1209] = 4'b0000;
	mem[1210] = 4'b0000;
	mem[1211] = 4'b0001;
	mem[1212] = 4'b0001;
	mem[1213] = 4'b0000;
	mem[1214] = 4'b0000;
	mem[1215] = 4'b0000;
	mem[1216] = 4'b0000;
	mem[1217] = 4'b0001;
	mem[1218] = 4'b0000;
	mem[1219] = 4'b0000;
	mem[1220] = 4'b0000;
	mem[1221] = 4'b0000;
	mem[1222] = 4'b0000;
	mem[1223] = 4'b1100;
	mem[1224] = 4'b1111;
	mem[1225] = 4'b1111;
	mem[1226] = 4'b1111;
	mem[1227] = 4'b1111;
	mem[1228] = 4'b1111;
	mem[1229] = 4'b1111;
	mem[1230] = 4'b1111;
	mem[1231] = 4'b1111;
	mem[1232] = 4'b1111;
	mem[1233] = 4'b1111;
	mem[1234] = 4'b1111;
	mem[1235] = 4'b1111;
	mem[1236] = 4'b1111;
	mem[1237] = 4'b1111;
	mem[1238] = 4'b1111;
	mem[1239] = 4'b1111;
	mem[1240] = 4'b0100;
	mem[1241] = 4'b0000;
	mem[1242] = 4'b0000;
	mem[1243] = 4'b0000;
	mem[1244] = 4'b0000;
	mem[1245] = 4'b0000;
	mem[1246] = 4'b0000;
	mem[1247] = 4'b0000;
	mem[1248] = 4'b0000;
	mem[1249] = 4'b0000;
	mem[1250] = 4'b0000;
	mem[1251] = 4'b0000;
	mem[1252] = 4'b0001;
	mem[1253] = 4'b0001;
	mem[1254] = 4'b0000;
	mem[1255] = 4'b0000;
	mem[1256] = 4'b0000;
	mem[1257] = 4'b1000;
	mem[1258] = 4'b1111;
	mem[1259] = 4'b1111;
	mem[1260] = 4'b1111;
	mem[1261] = 4'b1111;
	mem[1262] = 4'b1110;
	mem[1263] = 4'b1111;
	mem[1264] = 4'b1111;
	mem[1265] = 4'b1111;
	mem[1266] = 4'b1111;
	mem[1267] = 4'b1111;
	mem[1268] = 4'b1111;
	mem[1269] = 4'b1111;
	mem[1270] = 4'b1111;
	mem[1271] = 4'b1111;
	mem[1272] = 4'b1111;
	mem[1273] = 4'b1111;
	mem[1274] = 4'b0011;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0111;
	mem[1284] = 4'b1100;
	mem[1285] = 4'b1101;
	mem[1286] = 4'b1110;
	mem[1287] = 4'b1110;
	mem[1288] = 4'b1110;
	mem[1289] = 4'b1110;
	mem[1290] = 4'b1110;
	mem[1291] = 4'b1101;
	mem[1292] = 4'b1100;
	mem[1293] = 4'b1100;
	mem[1294] = 4'b1100;
	mem[1295] = 4'b1100;
	mem[1296] = 4'b1100;
	mem[1297] = 4'b1100;
	mem[1298] = 4'b1100;
	mem[1299] = 4'b1100;
	mem[1300] = 4'b0011;
	mem[1301] = 4'b0000;
	mem[1302] = 4'b0000;
	mem[1303] = 4'b0000;
	mem[1304] = 4'b0000;
	mem[1305] = 4'b0000;
	mem[1306] = 4'b0000;
	mem[1307] = 4'b0000;
	mem[1308] = 4'b0000;
	mem[1309] = 4'b0000;
	mem[1310] = 4'b0000;
	mem[1311] = 4'b0000;
	mem[1312] = 4'b0000;
	mem[1313] = 4'b0000;
	mem[1314] = 4'b0000;
	mem[1315] = 4'b0000;
	mem[1316] = 4'b0000;
	mem[1317] = 4'b1100;
	mem[1318] = 4'b1111;
	mem[1319] = 4'b1111;
	mem[1320] = 4'b1111;
	mem[1321] = 4'b1111;
	mem[1322] = 4'b1111;
	mem[1323] = 4'b1111;
	mem[1324] = 4'b1111;
	mem[1325] = 4'b1111;
	mem[1326] = 4'b1111;
	mem[1327] = 4'b1111;
	mem[1328] = 4'b1111;
	mem[1329] = 4'b1111;
	mem[1330] = 4'b1101;
	mem[1331] = 4'b1101;
	mem[1332] = 4'b1101;
	mem[1333] = 4'b1101;
	mem[1334] = 4'b0101;
	mem[1335] = 4'b0000;
	mem[1336] = 4'b0000;
	mem[1337] = 4'b0001;
	mem[1338] = 4'b0001;
	mem[1339] = 4'b0000;
	mem[1340] = 4'b0000;
	mem[1341] = 4'b0000;
	mem[1342] = 4'b0000;
	mem[1343] = 4'b0000;
	mem[1344] = 4'b0000;
	mem[1345] = 4'b0001;
	mem[1346] = 4'b0000;
	mem[1347] = 4'b0000;
	mem[1348] = 4'b0000;
	mem[1349] = 4'b0000;
	mem[1350] = 4'b0000;
	mem[1351] = 4'b1100;
	mem[1352] = 4'b1111;
	mem[1353] = 4'b1111;
	mem[1354] = 4'b1111;
	mem[1355] = 4'b1111;
	mem[1356] = 4'b1111;
	mem[1357] = 4'b1111;
	mem[1358] = 4'b1111;
	mem[1359] = 4'b1111;
	mem[1360] = 4'b1111;
	mem[1361] = 4'b1111;
	mem[1362] = 4'b1111;
	mem[1363] = 4'b1111;
	mem[1364] = 4'b1111;
	mem[1365] = 4'b1111;
	mem[1366] = 4'b1111;
	mem[1367] = 4'b1111;
	mem[1368] = 4'b0100;
	mem[1369] = 4'b0000;
	mem[1370] = 4'b0000;
	mem[1371] = 4'b0000;
	mem[1372] = 4'b0000;
	mem[1373] = 4'b0000;
	mem[1374] = 4'b0000;
	mem[1375] = 4'b0000;
	mem[1376] = 4'b0000;
	mem[1377] = 4'b0000;
	mem[1378] = 4'b0000;
	mem[1379] = 4'b0000;
	mem[1380] = 4'b0001;
	mem[1381] = 4'b0000;
	mem[1382] = 4'b0000;
	mem[1383] = 4'b0000;
	mem[1384] = 4'b0001;
	mem[1385] = 4'b1000;
	mem[1386] = 4'b1101;
	mem[1387] = 4'b1111;
	mem[1388] = 4'b1111;
	mem[1389] = 4'b1111;
	mem[1390] = 4'b1111;
	mem[1391] = 4'b1111;
	mem[1392] = 4'b1111;
	mem[1393] = 4'b1111;
	mem[1394] = 4'b1111;
	mem[1395] = 4'b1111;
	mem[1396] = 4'b1111;
	mem[1397] = 4'b1111;
	mem[1398] = 4'b1111;
	mem[1399] = 4'b1111;
	mem[1400] = 4'b1111;
	mem[1401] = 4'b1111;
	mem[1402] = 4'b0011;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0111;
	mem[1412] = 4'b1100;
	mem[1413] = 4'b1101;
	mem[1414] = 4'b1110;
	mem[1415] = 4'b1110;
	mem[1416] = 4'b1110;
	mem[1417] = 4'b1101;
	mem[1418] = 4'b1100;
	mem[1419] = 4'b1100;
	mem[1420] = 4'b1100;
	mem[1421] = 4'b1100;
	mem[1422] = 4'b1100;
	mem[1423] = 4'b1100;
	mem[1424] = 4'b1100;
	mem[1425] = 4'b1100;
	mem[1426] = 4'b1100;
	mem[1427] = 4'b1100;
	mem[1428] = 4'b0011;
	mem[1429] = 4'b0000;
	mem[1430] = 4'b0000;
	mem[1431] = 4'b0000;
	mem[1432] = 4'b0000;
	mem[1433] = 4'b0000;
	mem[1434] = 4'b0000;
	mem[1435] = 4'b0000;
	mem[1436] = 4'b0000;
	mem[1437] = 4'b0000;
	mem[1438] = 4'b0000;
	mem[1439] = 4'b0000;
	mem[1440] = 4'b0000;
	mem[1441] = 4'b0000;
	mem[1442] = 4'b0000;
	mem[1443] = 4'b0000;
	mem[1444] = 4'b0000;
	mem[1445] = 4'b1100;
	mem[1446] = 4'b1111;
	mem[1447] = 4'b1111;
	mem[1448] = 4'b1111;
	mem[1449] = 4'b1111;
	mem[1450] = 4'b1111;
	mem[1451] = 4'b1111;
	mem[1452] = 4'b1111;
	mem[1453] = 4'b1111;
	mem[1454] = 4'b1111;
	mem[1455] = 4'b1111;
	mem[1456] = 4'b1111;
	mem[1457] = 4'b1111;
	mem[1458] = 4'b1111;
	mem[1459] = 4'b1110;
	mem[1460] = 4'b1101;
	mem[1461] = 4'b1101;
	mem[1462] = 4'b0101;
	mem[1463] = 4'b0001;
	mem[1464] = 4'b0001;
	mem[1465] = 4'b0000;
	mem[1466] = 4'b0000;
	mem[1467] = 4'b0000;
	mem[1468] = 4'b0000;
	mem[1469] = 4'b0000;
	mem[1470] = 4'b0000;
	mem[1471] = 4'b0000;
	mem[1472] = 4'b0001;
	mem[1473] = 4'b0001;
	mem[1474] = 4'b0000;
	mem[1475] = 4'b0000;
	mem[1476] = 4'b0000;
	mem[1477] = 4'b0000;
	mem[1478] = 4'b0000;
	mem[1479] = 4'b1100;
	mem[1480] = 4'b1111;
	mem[1481] = 4'b1111;
	mem[1482] = 4'b1111;
	mem[1483] = 4'b1111;
	mem[1484] = 4'b1111;
	mem[1485] = 4'b1111;
	mem[1486] = 4'b1111;
	mem[1487] = 4'b1111;
	mem[1488] = 4'b1111;
	mem[1489] = 4'b1111;
	mem[1490] = 4'b1111;
	mem[1491] = 4'b1111;
	mem[1492] = 4'b1111;
	mem[1493] = 4'b1111;
	mem[1494] = 4'b1111;
	mem[1495] = 4'b1111;
	mem[1496] = 4'b0100;
	mem[1497] = 4'b0000;
	mem[1498] = 4'b0000;
	mem[1499] = 4'b0000;
	mem[1500] = 4'b0000;
	mem[1501] = 4'b0000;
	mem[1502] = 4'b0000;
	mem[1503] = 4'b0000;
	mem[1504] = 4'b0000;
	mem[1505] = 4'b0000;
	mem[1506] = 4'b0000;
	mem[1507] = 4'b0000;
	mem[1508] = 4'b0001;
	mem[1509] = 4'b0000;
	mem[1510] = 4'b0000;
	mem[1511] = 4'b0001;
	mem[1512] = 4'b0001;
	mem[1513] = 4'b1001;
	mem[1514] = 4'b1101;
	mem[1515] = 4'b1101;
	mem[1516] = 4'b1110;
	mem[1517] = 4'b1111;
	mem[1518] = 4'b1111;
	mem[1519] = 4'b1111;
	mem[1520] = 4'b1111;
	mem[1521] = 4'b1111;
	mem[1522] = 4'b1111;
	mem[1523] = 4'b1111;
	mem[1524] = 4'b1111;
	mem[1525] = 4'b1111;
	mem[1526] = 4'b1111;
	mem[1527] = 4'b1111;
	mem[1528] = 4'b1111;
	mem[1529] = 4'b1111;
	mem[1530] = 4'b0011;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b1001;
	mem[1540] = 4'b1111;
	mem[1541] = 4'b1111;
	mem[1542] = 4'b1111;
	mem[1543] = 4'b1111;
	mem[1544] = 4'b1111;
	mem[1545] = 4'b1111;
	mem[1546] = 4'b1111;
	mem[1547] = 4'b1111;
	mem[1548] = 4'b1111;
	mem[1549] = 4'b1111;
	mem[1550] = 4'b1111;
	mem[1551] = 4'b1111;
	mem[1552] = 4'b1111;
	mem[1553] = 4'b1111;
	mem[1554] = 4'b1111;
	mem[1555] = 4'b1111;
	mem[1556] = 4'b0011;
	mem[1557] = 4'b0000;
	mem[1558] = 4'b0000;
	mem[1559] = 4'b0000;
	mem[1560] = 4'b0000;
	mem[1561] = 4'b0000;
	mem[1562] = 4'b0000;
	mem[1563] = 4'b0000;
	mem[1564] = 4'b0000;
	mem[1565] = 4'b0000;
	mem[1566] = 4'b0000;
	mem[1567] = 4'b0000;
	mem[1568] = 4'b0000;
	mem[1569] = 4'b0000;
	mem[1570] = 4'b0000;
	mem[1571] = 4'b0000;
	mem[1572] = 4'b0000;
	mem[1573] = 4'b1100;
	mem[1574] = 4'b1111;
	mem[1575] = 4'b1111;
	mem[1576] = 4'b1111;
	mem[1577] = 4'b1111;
	mem[1578] = 4'b1111;
	mem[1579] = 4'b1110;
	mem[1580] = 4'b1101;
	mem[1581] = 4'b1110;
	mem[1582] = 4'b1110;
	mem[1583] = 4'b1111;
	mem[1584] = 4'b1111;
	mem[1585] = 4'b1111;
	mem[1586] = 4'b1111;
	mem[1587] = 4'b1111;
	mem[1588] = 4'b1111;
	mem[1589] = 4'b1111;
	mem[1590] = 4'b0110;
	mem[1591] = 4'b0000;
	mem[1592] = 4'b0000;
	mem[1593] = 4'b0000;
	mem[1594] = 4'b0000;
	mem[1595] = 4'b0000;
	mem[1596] = 4'b0000;
	mem[1597] = 4'b0000;
	mem[1598] = 4'b0000;
	mem[1599] = 4'b0000;
	mem[1600] = 4'b0001;
	mem[1601] = 4'b0000;
	mem[1602] = 4'b0000;
	mem[1603] = 4'b0000;
	mem[1604] = 4'b0000;
	mem[1605] = 4'b0000;
	mem[1606] = 4'b0000;
	mem[1607] = 4'b1100;
	mem[1608] = 4'b1111;
	mem[1609] = 4'b1111;
	mem[1610] = 4'b1111;
	mem[1611] = 4'b1111;
	mem[1612] = 4'b1111;
	mem[1613] = 4'b1111;
	mem[1614] = 4'b1111;
	mem[1615] = 4'b1111;
	mem[1616] = 4'b1111;
	mem[1617] = 4'b1111;
	mem[1618] = 4'b1111;
	mem[1619] = 4'b1111;
	mem[1620] = 4'b1111;
	mem[1621] = 4'b1111;
	mem[1622] = 4'b1111;
	mem[1623] = 4'b1111;
	mem[1624] = 4'b0100;
	mem[1625] = 4'b0000;
	mem[1626] = 4'b0000;
	mem[1627] = 4'b0000;
	mem[1628] = 4'b0000;
	mem[1629] = 4'b0000;
	mem[1630] = 4'b0000;
	mem[1631] = 4'b0000;
	mem[1632] = 4'b0000;
	mem[1633] = 4'b0000;
	mem[1634] = 4'b0000;
	mem[1635] = 4'b0001;
	mem[1636] = 4'b0000;
	mem[1637] = 4'b0000;
	mem[1638] = 4'b0001;
	mem[1639] = 4'b0001;
	mem[1640] = 4'b0000;
	mem[1641] = 4'b0111;
	mem[1642] = 4'b1011;
	mem[1643] = 4'b1100;
	mem[1644] = 4'b1101;
	mem[1645] = 4'b1101;
	mem[1646] = 4'b1101;
	mem[1647] = 4'b1101;
	mem[1648] = 4'b1101;
	mem[1649] = 4'b1101;
	mem[1650] = 4'b1101;
	mem[1651] = 4'b1101;
	mem[1652] = 4'b1101;
	mem[1653] = 4'b1101;
	mem[1654] = 4'b1101;
	mem[1655] = 4'b1101;
	mem[1656] = 4'b1101;
	mem[1657] = 4'b1100;
	mem[1658] = 4'b0011;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b1001;
	mem[1668] = 4'b1111;
	mem[1669] = 4'b1111;
	mem[1670] = 4'b1111;
	mem[1671] = 4'b1111;
	mem[1672] = 4'b1111;
	mem[1673] = 4'b1111;
	mem[1674] = 4'b1111;
	mem[1675] = 4'b1111;
	mem[1676] = 4'b1111;
	mem[1677] = 4'b1111;
	mem[1678] = 4'b1111;
	mem[1679] = 4'b1111;
	mem[1680] = 4'b1111;
	mem[1681] = 4'b1111;
	mem[1682] = 4'b1111;
	mem[1683] = 4'b1111;
	mem[1684] = 4'b0100;
	mem[1685] = 4'b0000;
	mem[1686] = 4'b0000;
	mem[1687] = 4'b0000;
	mem[1688] = 4'b0000;
	mem[1689] = 4'b0000;
	mem[1690] = 4'b0000;
	mem[1691] = 4'b0000;
	mem[1692] = 4'b0000;
	mem[1693] = 4'b0000;
	mem[1694] = 4'b0000;
	mem[1695] = 4'b0000;
	mem[1696] = 4'b0000;
	mem[1697] = 4'b0000;
	mem[1698] = 4'b0000;
	mem[1699] = 4'b0000;
	mem[1700] = 4'b0000;
	mem[1701] = 4'b1100;
	mem[1702] = 4'b1111;
	mem[1703] = 4'b1111;
	mem[1704] = 4'b1111;
	mem[1705] = 4'b1110;
	mem[1706] = 4'b1101;
	mem[1707] = 4'b1101;
	mem[1708] = 4'b1101;
	mem[1709] = 4'b1101;
	mem[1710] = 4'b1101;
	mem[1711] = 4'b1101;
	mem[1712] = 4'b1111;
	mem[1713] = 4'b1111;
	mem[1714] = 4'b1111;
	mem[1715] = 4'b1111;
	mem[1716] = 4'b1111;
	mem[1717] = 4'b1111;
	mem[1718] = 4'b0110;
	mem[1719] = 4'b0000;
	mem[1720] = 4'b0000;
	mem[1721] = 4'b0000;
	mem[1722] = 4'b0000;
	mem[1723] = 4'b0000;
	mem[1724] = 4'b0000;
	mem[1725] = 4'b0000;
	mem[1726] = 4'b0000;
	mem[1727] = 4'b0001;
	mem[1728] = 4'b0001;
	mem[1729] = 4'b0000;
	mem[1730] = 4'b0000;
	mem[1731] = 4'b0000;
	mem[1732] = 4'b0000;
	mem[1733] = 4'b0000;
	mem[1734] = 4'b0000;
	mem[1735] = 4'b1100;
	mem[1736] = 4'b1111;
	mem[1737] = 4'b1111;
	mem[1738] = 4'b1111;
	mem[1739] = 4'b1111;
	mem[1740] = 4'b1111;
	mem[1741] = 4'b1111;
	mem[1742] = 4'b1111;
	mem[1743] = 4'b1111;
	mem[1744] = 4'b1111;
	mem[1745] = 4'b1111;
	mem[1746] = 4'b1111;
	mem[1747] = 4'b1111;
	mem[1748] = 4'b1111;
	mem[1749] = 4'b1111;
	mem[1750] = 4'b1111;
	mem[1751] = 4'b1111;
	mem[1752] = 4'b0100;
	mem[1753] = 4'b0000;
	mem[1754] = 4'b0000;
	mem[1755] = 4'b0000;
	mem[1756] = 4'b0000;
	mem[1757] = 4'b0000;
	mem[1758] = 4'b0000;
	mem[1759] = 4'b0000;
	mem[1760] = 4'b0000;
	mem[1761] = 4'b0000;
	mem[1762] = 4'b0000;
	mem[1763] = 4'b0000;
	mem[1764] = 4'b0000;
	mem[1765] = 4'b0000;
	mem[1766] = 4'b0000;
	mem[1767] = 4'b0000;
	mem[1768] = 4'b0000;
	mem[1769] = 4'b0111;
	mem[1770] = 4'b1100;
	mem[1771] = 4'b1100;
	mem[1772] = 4'b1100;
	mem[1773] = 4'b1100;
	mem[1774] = 4'b1100;
	mem[1775] = 4'b1100;
	mem[1776] = 4'b1100;
	mem[1777] = 4'b1100;
	mem[1778] = 4'b1100;
	mem[1779] = 4'b1100;
	mem[1780] = 4'b1100;
	mem[1781] = 4'b1100;
	mem[1782] = 4'b1100;
	mem[1783] = 4'b1100;
	mem[1784] = 4'b1100;
	mem[1785] = 4'b1100;
	mem[1786] = 4'b0010;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b1001;
	mem[1796] = 4'b1111;
	mem[1797] = 4'b1111;
	mem[1798] = 4'b1111;
	mem[1799] = 4'b1111;
	mem[1800] = 4'b1111;
	mem[1801] = 4'b1111;
	mem[1802] = 4'b1111;
	mem[1803] = 4'b1111;
	mem[1804] = 4'b1111;
	mem[1805] = 4'b1111;
	mem[1806] = 4'b1111;
	mem[1807] = 4'b1111;
	mem[1808] = 4'b1111;
	mem[1809] = 4'b1111;
	mem[1810] = 4'b1111;
	mem[1811] = 4'b1111;
	mem[1812] = 4'b0100;
	mem[1813] = 4'b0000;
	mem[1814] = 4'b0000;
	mem[1815] = 4'b0000;
	mem[1816] = 4'b0000;
	mem[1817] = 4'b0000;
	mem[1818] = 4'b0000;
	mem[1819] = 4'b0000;
	mem[1820] = 4'b0000;
	mem[1821] = 4'b0000;
	mem[1822] = 4'b0000;
	mem[1823] = 4'b0000;
	mem[1824] = 4'b0000;
	mem[1825] = 4'b0000;
	mem[1826] = 4'b0000;
	mem[1827] = 4'b0000;
	mem[1828] = 4'b0000;
	mem[1829] = 4'b1100;
	mem[1830] = 4'b1111;
	mem[1831] = 4'b1111;
	mem[1832] = 4'b1110;
	mem[1833] = 4'b1101;
	mem[1834] = 4'b1101;
	mem[1835] = 4'b1101;
	mem[1836] = 4'b1101;
	mem[1837] = 4'b1101;
	mem[1838] = 4'b1101;
	mem[1839] = 4'b1101;
	mem[1840] = 4'b1101;
	mem[1841] = 4'b1111;
	mem[1842] = 4'b1111;
	mem[1843] = 4'b1111;
	mem[1844] = 4'b1111;
	mem[1845] = 4'b1111;
	mem[1846] = 4'b0110;
	mem[1847] = 4'b0000;
	mem[1848] = 4'b0000;
	mem[1849] = 4'b0000;
	mem[1850] = 4'b0000;
	mem[1851] = 4'b0000;
	mem[1852] = 4'b0000;
	mem[1853] = 4'b0000;
	mem[1854] = 4'b0001;
	mem[1855] = 4'b0001;
	mem[1856] = 4'b0000;
	mem[1857] = 4'b0000;
	mem[1858] = 4'b0000;
	mem[1859] = 4'b0000;
	mem[1860] = 4'b0000;
	mem[1861] = 4'b0000;
	mem[1862] = 4'b0000;
	mem[1863] = 4'b1100;
	mem[1864] = 4'b1111;
	mem[1865] = 4'b1111;
	mem[1866] = 4'b1111;
	mem[1867] = 4'b1111;
	mem[1868] = 4'b1111;
	mem[1869] = 4'b1111;
	mem[1870] = 4'b1111;
	mem[1871] = 4'b1111;
	mem[1872] = 4'b1111;
	mem[1873] = 4'b1111;
	mem[1874] = 4'b1111;
	mem[1875] = 4'b1111;
	mem[1876] = 4'b1111;
	mem[1877] = 4'b1111;
	mem[1878] = 4'b1111;
	mem[1879] = 4'b1111;
	mem[1880] = 4'b0011;
	mem[1881] = 4'b0000;
	mem[1882] = 4'b0000;
	mem[1883] = 4'b0000;
	mem[1884] = 4'b0000;
	mem[1885] = 4'b0000;
	mem[1886] = 4'b0000;
	mem[1887] = 4'b0000;
	mem[1888] = 4'b0000;
	mem[1889] = 4'b0000;
	mem[1890] = 4'b0000;
	mem[1891] = 4'b0000;
	mem[1892] = 4'b0000;
	mem[1893] = 4'b0000;
	mem[1894] = 4'b0000;
	mem[1895] = 4'b0000;
	mem[1896] = 4'b0000;
	mem[1897] = 4'b0111;
	mem[1898] = 4'b1101;
	mem[1899] = 4'b1100;
	mem[1900] = 4'b1100;
	mem[1901] = 4'b1100;
	mem[1902] = 4'b1100;
	mem[1903] = 4'b1100;
	mem[1904] = 4'b1100;
	mem[1905] = 4'b1100;
	mem[1906] = 4'b1100;
	mem[1907] = 4'b1100;
	mem[1908] = 4'b1100;
	mem[1909] = 4'b1100;
	mem[1910] = 4'b1100;
	mem[1911] = 4'b1100;
	mem[1912] = 4'b1100;
	mem[1913] = 4'b1100;
	mem[1914] = 4'b0010;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b1001;
	mem[1924] = 4'b1111;
	mem[1925] = 4'b1111;
	mem[1926] = 4'b1111;
	mem[1927] = 4'b1111;
	mem[1928] = 4'b1111;
	mem[1929] = 4'b1111;
	mem[1930] = 4'b1111;
	mem[1931] = 4'b1111;
	mem[1932] = 4'b1111;
	mem[1933] = 4'b1111;
	mem[1934] = 4'b1111;
	mem[1935] = 4'b1111;
	mem[1936] = 4'b1111;
	mem[1937] = 4'b1111;
	mem[1938] = 4'b1111;
	mem[1939] = 4'b1111;
	mem[1940] = 4'b0100;
	mem[1941] = 4'b0000;
	mem[1942] = 4'b0000;
	mem[1943] = 4'b0000;
	mem[1944] = 4'b0000;
	mem[1945] = 4'b0000;
	mem[1946] = 4'b0000;
	mem[1947] = 4'b0000;
	mem[1948] = 4'b0000;
	mem[1949] = 4'b0000;
	mem[1950] = 4'b0000;
	mem[1951] = 4'b0000;
	mem[1952] = 4'b0000;
	mem[1953] = 4'b0000;
	mem[1954] = 4'b0000;
	mem[1955] = 4'b0000;
	mem[1956] = 4'b0000;
	mem[1957] = 4'b1100;
	mem[1958] = 4'b1111;
	mem[1959] = 4'b1111;
	mem[1960] = 4'b1101;
	mem[1961] = 4'b1101;
	mem[1962] = 4'b1101;
	mem[1963] = 4'b1101;
	mem[1964] = 4'b1101;
	mem[1965] = 4'b1101;
	mem[1966] = 4'b1101;
	mem[1967] = 4'b1101;
	mem[1968] = 4'b1101;
	mem[1969] = 4'b1101;
	mem[1970] = 4'b1111;
	mem[1971] = 4'b1111;
	mem[1972] = 4'b1111;
	mem[1973] = 4'b1111;
	mem[1974] = 4'b0101;
	mem[1975] = 4'b0000;
	mem[1976] = 4'b0000;
	mem[1977] = 4'b0000;
	mem[1978] = 4'b0000;
	mem[1979] = 4'b0000;
	mem[1980] = 4'b0000;
	mem[1981] = 4'b0001;
	mem[1982] = 4'b0001;
	mem[1983] = 4'b0000;
	mem[1984] = 4'b0000;
	mem[1985] = 4'b0000;
	mem[1986] = 4'b0000;
	mem[1987] = 4'b0000;
	mem[1988] = 4'b0000;
	mem[1989] = 4'b0000;
	mem[1990] = 4'b0000;
	mem[1991] = 4'b1100;
	mem[1992] = 4'b1111;
	mem[1993] = 4'b1111;
	mem[1994] = 4'b1111;
	mem[1995] = 4'b1111;
	mem[1996] = 4'b1111;
	mem[1997] = 4'b1111;
	mem[1998] = 4'b1111;
	mem[1999] = 4'b1111;
	mem[2000] = 4'b1111;
	mem[2001] = 4'b1111;
	mem[2002] = 4'b1111;
	mem[2003] = 4'b1111;
	mem[2004] = 4'b1111;
	mem[2005] = 4'b1111;
	mem[2006] = 4'b1111;
	mem[2007] = 4'b1111;
	mem[2008] = 4'b0100;
	mem[2009] = 4'b0000;
	mem[2010] = 4'b0000;
	mem[2011] = 4'b0000;
	mem[2012] = 4'b0000;
	mem[2013] = 4'b0000;
	mem[2014] = 4'b0000;
	mem[2015] = 4'b0000;
	mem[2016] = 4'b0000;
	mem[2017] = 4'b0000;
	mem[2018] = 4'b0000;
	mem[2019] = 4'b0000;
	mem[2020] = 4'b0000;
	mem[2021] = 4'b0000;
	mem[2022] = 4'b0000;
	mem[2023] = 4'b0000;
	mem[2024] = 4'b0001;
	mem[2025] = 4'b1000;
	mem[2026] = 4'b1100;
	mem[2027] = 4'b1100;
	mem[2028] = 4'b1100;
	mem[2029] = 4'b1100;
	mem[2030] = 4'b1100;
	mem[2031] = 4'b1100;
	mem[2032] = 4'b1100;
	mem[2033] = 4'b1100;
	mem[2034] = 4'b1100;
	mem[2035] = 4'b1100;
	mem[2036] = 4'b1100;
	mem[2037] = 4'b1100;
	mem[2038] = 4'b1100;
	mem[2039] = 4'b1100;
	mem[2040] = 4'b1100;
	mem[2041] = 4'b1100;
	mem[2042] = 4'b0010;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b1001;
	mem[2052] = 4'b1111;
	mem[2053] = 4'b1111;
	mem[2054] = 4'b1111;
	mem[2055] = 4'b1111;
	mem[2056] = 4'b1111;
	mem[2057] = 4'b1111;
	mem[2058] = 4'b1111;
	mem[2059] = 4'b1111;
	mem[2060] = 4'b1111;
	mem[2061] = 4'b1111;
	mem[2062] = 4'b1111;
	mem[2063] = 4'b1111;
	mem[2064] = 4'b1111;
	mem[2065] = 4'b1111;
	mem[2066] = 4'b1111;
	mem[2067] = 4'b1111;
	mem[2068] = 4'b0100;
	mem[2069] = 4'b0000;
	mem[2070] = 4'b0000;
	mem[2071] = 4'b0000;
	mem[2072] = 4'b0000;
	mem[2073] = 4'b0000;
	mem[2074] = 4'b0000;
	mem[2075] = 4'b0000;
	mem[2076] = 4'b0000;
	mem[2077] = 4'b0000;
	mem[2078] = 4'b0000;
	mem[2079] = 4'b0000;
	mem[2080] = 4'b0000;
	mem[2081] = 4'b0000;
	mem[2082] = 4'b0000;
	mem[2083] = 4'b0000;
	mem[2084] = 4'b0000;
	mem[2085] = 4'b1100;
	mem[2086] = 4'b1111;
	mem[2087] = 4'b1111;
	mem[2088] = 4'b1101;
	mem[2089] = 4'b1101;
	mem[2090] = 4'b1110;
	mem[2091] = 4'b1111;
	mem[2092] = 4'b1111;
	mem[2093] = 4'b1111;
	mem[2094] = 4'b1101;
	mem[2095] = 4'b1101;
	mem[2096] = 4'b1101;
	mem[2097] = 4'b1101;
	mem[2098] = 4'b1101;
	mem[2099] = 4'b1111;
	mem[2100] = 4'b1111;
	mem[2101] = 4'b1111;
	mem[2102] = 4'b0110;
	mem[2103] = 4'b0001;
	mem[2104] = 4'b0001;
	mem[2105] = 4'b0000;
	mem[2106] = 4'b0001;
	mem[2107] = 4'b0001;
	mem[2108] = 4'b0001;
	mem[2109] = 4'b0000;
	mem[2110] = 4'b0000;
	mem[2111] = 4'b0000;
	mem[2112] = 4'b0000;
	mem[2113] = 4'b0000;
	mem[2114] = 4'b0000;
	mem[2115] = 4'b0000;
	mem[2116] = 4'b0000;
	mem[2117] = 4'b0000;
	mem[2118] = 4'b0000;
	mem[2119] = 4'b1100;
	mem[2120] = 4'b1111;
	mem[2121] = 4'b1111;
	mem[2122] = 4'b1111;
	mem[2123] = 4'b1111;
	mem[2124] = 4'b1111;
	mem[2125] = 4'b1111;
	mem[2126] = 4'b1111;
	mem[2127] = 4'b1111;
	mem[2128] = 4'b1111;
	mem[2129] = 4'b1111;
	mem[2130] = 4'b1111;
	mem[2131] = 4'b1111;
	mem[2132] = 4'b1111;
	mem[2133] = 4'b1111;
	mem[2134] = 4'b1111;
	mem[2135] = 4'b1111;
	mem[2136] = 4'b0100;
	mem[2137] = 4'b0000;
	mem[2138] = 4'b0000;
	mem[2139] = 4'b0000;
	mem[2140] = 4'b0000;
	mem[2141] = 4'b0000;
	mem[2142] = 4'b0000;
	mem[2143] = 4'b0000;
	mem[2144] = 4'b0000;
	mem[2145] = 4'b0000;
	mem[2146] = 4'b0000;
	mem[2147] = 4'b0000;
	mem[2148] = 4'b0000;
	mem[2149] = 4'b0000;
	mem[2150] = 4'b0000;
	mem[2151] = 4'b0001;
	mem[2152] = 4'b0001;
	mem[2153] = 4'b1000;
	mem[2154] = 4'b1100;
	mem[2155] = 4'b1100;
	mem[2156] = 4'b1100;
	mem[2157] = 4'b1100;
	mem[2158] = 4'b1100;
	mem[2159] = 4'b1100;
	mem[2160] = 4'b1100;
	mem[2161] = 4'b1100;
	mem[2162] = 4'b1100;
	mem[2163] = 4'b1100;
	mem[2164] = 4'b1100;
	mem[2165] = 4'b1100;
	mem[2166] = 4'b1100;
	mem[2167] = 4'b1100;
	mem[2168] = 4'b1100;
	mem[2169] = 4'b1100;
	mem[2170] = 4'b0010;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b1001;
	mem[2180] = 4'b1111;
	mem[2181] = 4'b1111;
	mem[2182] = 4'b1111;
	mem[2183] = 4'b1111;
	mem[2184] = 4'b1111;
	mem[2185] = 4'b1111;
	mem[2186] = 4'b1111;
	mem[2187] = 4'b1111;
	mem[2188] = 4'b1111;
	mem[2189] = 4'b1111;
	mem[2190] = 4'b1111;
	mem[2191] = 4'b1111;
	mem[2192] = 4'b1111;
	mem[2193] = 4'b1111;
	mem[2194] = 4'b1111;
	mem[2195] = 4'b1111;
	mem[2196] = 4'b0100;
	mem[2197] = 4'b0000;
	mem[2198] = 4'b0000;
	mem[2199] = 4'b0000;
	mem[2200] = 4'b0000;
	mem[2201] = 4'b0000;
	mem[2202] = 4'b0000;
	mem[2203] = 4'b0000;
	mem[2204] = 4'b0000;
	mem[2205] = 4'b0000;
	mem[2206] = 4'b0000;
	mem[2207] = 4'b0000;
	mem[2208] = 4'b0000;
	mem[2209] = 4'b0000;
	mem[2210] = 4'b0000;
	mem[2211] = 4'b0000;
	mem[2212] = 4'b0000;
	mem[2213] = 4'b1011;
	mem[2214] = 4'b1111;
	mem[2215] = 4'b1111;
	mem[2216] = 4'b1101;
	mem[2217] = 4'b1110;
	mem[2218] = 4'b1111;
	mem[2219] = 4'b1111;
	mem[2220] = 4'b1111;
	mem[2221] = 4'b1111;
	mem[2222] = 4'b1111;
	mem[2223] = 4'b1101;
	mem[2224] = 4'b1101;
	mem[2225] = 4'b1101;
	mem[2226] = 4'b1101;
	mem[2227] = 4'b1101;
	mem[2228] = 4'b1111;
	mem[2229] = 4'b1111;
	mem[2230] = 4'b0110;
	mem[2231] = 4'b0000;
	mem[2232] = 4'b0000;
	mem[2233] = 4'b0000;
	mem[2234] = 4'b0000;
	mem[2235] = 4'b0000;
	mem[2236] = 4'b0000;
	mem[2237] = 4'b0000;
	mem[2238] = 4'b0000;
	mem[2239] = 4'b0000;
	mem[2240] = 4'b0000;
	mem[2241] = 4'b0000;
	mem[2242] = 4'b0000;
	mem[2243] = 4'b0000;
	mem[2244] = 4'b0000;
	mem[2245] = 4'b0000;
	mem[2246] = 4'b0000;
	mem[2247] = 4'b1100;
	mem[2248] = 4'b1111;
	mem[2249] = 4'b1111;
	mem[2250] = 4'b1111;
	mem[2251] = 4'b1111;
	mem[2252] = 4'b1111;
	mem[2253] = 4'b1111;
	mem[2254] = 4'b1111;
	mem[2255] = 4'b1111;
	mem[2256] = 4'b1111;
	mem[2257] = 4'b1111;
	mem[2258] = 4'b1111;
	mem[2259] = 4'b1111;
	mem[2260] = 4'b1111;
	mem[2261] = 4'b1111;
	mem[2262] = 4'b1111;
	mem[2263] = 4'b1111;
	mem[2264] = 4'b0100;
	mem[2265] = 4'b0000;
	mem[2266] = 4'b0000;
	mem[2267] = 4'b0000;
	mem[2268] = 4'b0000;
	mem[2269] = 4'b0000;
	mem[2270] = 4'b0000;
	mem[2271] = 4'b0000;
	mem[2272] = 4'b0000;
	mem[2273] = 4'b0000;
	mem[2274] = 4'b0000;
	mem[2275] = 4'b0000;
	mem[2276] = 4'b0000;
	mem[2277] = 4'b0000;
	mem[2278] = 4'b0000;
	mem[2279] = 4'b0000;
	mem[2280] = 4'b0000;
	mem[2281] = 4'b1000;
	mem[2282] = 4'b1100;
	mem[2283] = 4'b1100;
	mem[2284] = 4'b1100;
	mem[2285] = 4'b1100;
	mem[2286] = 4'b1100;
	mem[2287] = 4'b1100;
	mem[2288] = 4'b1100;
	mem[2289] = 4'b1100;
	mem[2290] = 4'b1100;
	mem[2291] = 4'b1100;
	mem[2292] = 4'b1100;
	mem[2293] = 4'b1100;
	mem[2294] = 4'b1100;
	mem[2295] = 4'b1100;
	mem[2296] = 4'b1100;
	mem[2297] = 4'b1100;
	mem[2298] = 4'b0010;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b1001;
	mem[2308] = 4'b1111;
	mem[2309] = 4'b1111;
	mem[2310] = 4'b1111;
	mem[2311] = 4'b1111;
	mem[2312] = 4'b1111;
	mem[2313] = 4'b1111;
	mem[2314] = 4'b1111;
	mem[2315] = 4'b1111;
	mem[2316] = 4'b1111;
	mem[2317] = 4'b1111;
	mem[2318] = 4'b1111;
	mem[2319] = 4'b1111;
	mem[2320] = 4'b1111;
	mem[2321] = 4'b1111;
	mem[2322] = 4'b1111;
	mem[2323] = 4'b1111;
	mem[2324] = 4'b0100;
	mem[2325] = 4'b0000;
	mem[2326] = 4'b0000;
	mem[2327] = 4'b0000;
	mem[2328] = 4'b0000;
	mem[2329] = 4'b0000;
	mem[2330] = 4'b0000;
	mem[2331] = 4'b0000;
	mem[2332] = 4'b0000;
	mem[2333] = 4'b0000;
	mem[2334] = 4'b0000;
	mem[2335] = 4'b0000;
	mem[2336] = 4'b0000;
	mem[2337] = 4'b0000;
	mem[2338] = 4'b0000;
	mem[2339] = 4'b0000;
	mem[2340] = 4'b0000;
	mem[2341] = 4'b1010;
	mem[2342] = 4'b1110;
	mem[2343] = 4'b1110;
	mem[2344] = 4'b1101;
	mem[2345] = 4'b1111;
	mem[2346] = 4'b1111;
	mem[2347] = 4'b1111;
	mem[2348] = 4'b1111;
	mem[2349] = 4'b1111;
	mem[2350] = 4'b1111;
	mem[2351] = 4'b1111;
	mem[2352] = 4'b1101;
	mem[2353] = 4'b1101;
	mem[2354] = 4'b1101;
	mem[2355] = 4'b1101;
	mem[2356] = 4'b1101;
	mem[2357] = 4'b1111;
	mem[2358] = 4'b0110;
	mem[2359] = 4'b0000;
	mem[2360] = 4'b0000;
	mem[2361] = 4'b0000;
	mem[2362] = 4'b0000;
	mem[2363] = 4'b0000;
	mem[2364] = 4'b0000;
	mem[2365] = 4'b0000;
	mem[2366] = 4'b0000;
	mem[2367] = 4'b0000;
	mem[2368] = 4'b0000;
	mem[2369] = 4'b0000;
	mem[2370] = 4'b0000;
	mem[2371] = 4'b0000;
	mem[2372] = 4'b0000;
	mem[2373] = 4'b0000;
	mem[2374] = 4'b0000;
	mem[2375] = 4'b1100;
	mem[2376] = 4'b1111;
	mem[2377] = 4'b1111;
	mem[2378] = 4'b1111;
	mem[2379] = 4'b1111;
	mem[2380] = 4'b1111;
	mem[2381] = 4'b1111;
	mem[2382] = 4'b1111;
	mem[2383] = 4'b1111;
	mem[2384] = 4'b1111;
	mem[2385] = 4'b1111;
	mem[2386] = 4'b1111;
	mem[2387] = 4'b1111;
	mem[2388] = 4'b1111;
	mem[2389] = 4'b1111;
	mem[2390] = 4'b1111;
	mem[2391] = 4'b1111;
	mem[2392] = 4'b0100;
	mem[2393] = 4'b0000;
	mem[2394] = 4'b0000;
	mem[2395] = 4'b0000;
	mem[2396] = 4'b0000;
	mem[2397] = 4'b0000;
	mem[2398] = 4'b0000;
	mem[2399] = 4'b0000;
	mem[2400] = 4'b0000;
	mem[2401] = 4'b0000;
	mem[2402] = 4'b0000;
	mem[2403] = 4'b0000;
	mem[2404] = 4'b0000;
	mem[2405] = 4'b0001;
	mem[2406] = 4'b0001;
	mem[2407] = 4'b0000;
	mem[2408] = 4'b0000;
	mem[2409] = 4'b1000;
	mem[2410] = 4'b1100;
	mem[2411] = 4'b1100;
	mem[2412] = 4'b1100;
	mem[2413] = 4'b1100;
	mem[2414] = 4'b1100;
	mem[2415] = 4'b1100;
	mem[2416] = 4'b1100;
	mem[2417] = 4'b1100;
	mem[2418] = 4'b1100;
	mem[2419] = 4'b1100;
	mem[2420] = 4'b1100;
	mem[2421] = 4'b1100;
	mem[2422] = 4'b1100;
	mem[2423] = 4'b1100;
	mem[2424] = 4'b1100;
	mem[2425] = 4'b1100;
	mem[2426] = 4'b0010;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b1001;
	mem[2436] = 4'b1111;
	mem[2437] = 4'b1111;
	mem[2438] = 4'b1111;
	mem[2439] = 4'b1111;
	mem[2440] = 4'b1111;
	mem[2441] = 4'b1111;
	mem[2442] = 4'b1111;
	mem[2443] = 4'b1111;
	mem[2444] = 4'b1111;
	mem[2445] = 4'b1111;
	mem[2446] = 4'b1111;
	mem[2447] = 4'b1111;
	mem[2448] = 4'b1111;
	mem[2449] = 4'b1111;
	mem[2450] = 4'b1111;
	mem[2451] = 4'b1111;
	mem[2452] = 4'b0100;
	mem[2453] = 4'b0000;
	mem[2454] = 4'b0000;
	mem[2455] = 4'b0000;
	mem[2456] = 4'b0000;
	mem[2457] = 4'b0000;
	mem[2458] = 4'b0000;
	mem[2459] = 4'b0000;
	mem[2460] = 4'b0000;
	mem[2461] = 4'b0000;
	mem[2462] = 4'b0000;
	mem[2463] = 4'b0000;
	mem[2464] = 4'b0000;
	mem[2465] = 4'b0000;
	mem[2466] = 4'b0000;
	mem[2467] = 4'b0000;
	mem[2468] = 4'b0000;
	mem[2469] = 4'b1010;
	mem[2470] = 4'b1101;
	mem[2471] = 4'b1101;
	mem[2472] = 4'b1101;
	mem[2473] = 4'b1111;
	mem[2474] = 4'b1111;
	mem[2475] = 4'b1111;
	mem[2476] = 4'b1111;
	mem[2477] = 4'b1111;
	mem[2478] = 4'b1111;
	mem[2479] = 4'b1111;
	mem[2480] = 4'b1111;
	mem[2481] = 4'b1101;
	mem[2482] = 4'b1101;
	mem[2483] = 4'b1101;
	mem[2484] = 4'b1101;
	mem[2485] = 4'b1101;
	mem[2486] = 4'b0110;
	mem[2487] = 4'b0000;
	mem[2488] = 4'b0000;
	mem[2489] = 4'b0000;
	mem[2490] = 4'b0000;
	mem[2491] = 4'b0000;
	mem[2492] = 4'b0000;
	mem[2493] = 4'b0000;
	mem[2494] = 4'b0000;
	mem[2495] = 4'b0000;
	mem[2496] = 4'b0000;
	mem[2497] = 4'b0000;
	mem[2498] = 4'b0000;
	mem[2499] = 4'b0000;
	mem[2500] = 4'b0000;
	mem[2501] = 4'b0000;
	mem[2502] = 4'b0000;
	mem[2503] = 4'b1100;
	mem[2504] = 4'b1111;
	mem[2505] = 4'b1111;
	mem[2506] = 4'b1111;
	mem[2507] = 4'b1111;
	mem[2508] = 4'b1111;
	mem[2509] = 4'b1111;
	mem[2510] = 4'b1111;
	mem[2511] = 4'b1111;
	mem[2512] = 4'b1111;
	mem[2513] = 4'b1111;
	mem[2514] = 4'b1111;
	mem[2515] = 4'b1111;
	mem[2516] = 4'b1111;
	mem[2517] = 4'b1111;
	mem[2518] = 4'b1111;
	mem[2519] = 4'b1111;
	mem[2520] = 4'b0100;
	mem[2521] = 4'b0000;
	mem[2522] = 4'b0000;
	mem[2523] = 4'b0000;
	mem[2524] = 4'b0000;
	mem[2525] = 4'b0000;
	mem[2526] = 4'b0000;
	mem[2527] = 4'b0000;
	mem[2528] = 4'b0000;
	mem[2529] = 4'b0000;
	mem[2530] = 4'b0000;
	mem[2531] = 4'b0000;
	mem[2532] = 4'b0001;
	mem[2533] = 4'b0001;
	mem[2534] = 4'b0000;
	mem[2535] = 4'b0000;
	mem[2536] = 4'b0000;
	mem[2537] = 4'b1000;
	mem[2538] = 4'b1100;
	mem[2539] = 4'b1100;
	mem[2540] = 4'b1100;
	mem[2541] = 4'b1100;
	mem[2542] = 4'b1100;
	mem[2543] = 4'b1100;
	mem[2544] = 4'b1100;
	mem[2545] = 4'b1100;
	mem[2546] = 4'b1100;
	mem[2547] = 4'b1100;
	mem[2548] = 4'b1100;
	mem[2549] = 4'b1100;
	mem[2550] = 4'b1100;
	mem[2551] = 4'b1100;
	mem[2552] = 4'b1100;
	mem[2553] = 4'b1100;
	mem[2554] = 4'b0010;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b1001;
	mem[2564] = 4'b1111;
	mem[2565] = 4'b1111;
	mem[2566] = 4'b1111;
	mem[2567] = 4'b1111;
	mem[2568] = 4'b1111;
	mem[2569] = 4'b1110;
	mem[2570] = 4'b1110;
	mem[2571] = 4'b1110;
	mem[2572] = 4'b1110;
	mem[2573] = 4'b1110;
	mem[2574] = 4'b1101;
	mem[2575] = 4'b1101;
	mem[2576] = 4'b1101;
	mem[2577] = 4'b1101;
	mem[2578] = 4'b1101;
	mem[2579] = 4'b1100;
	mem[2580] = 4'b1011;
	mem[2581] = 4'b1010;
	mem[2582] = 4'b1010;
	mem[2583] = 4'b1010;
	mem[2584] = 4'b1001;
	mem[2585] = 4'b1001;
	mem[2586] = 4'b1001;
	mem[2587] = 4'b1001;
	mem[2588] = 4'b1001;
	mem[2589] = 4'b1000;
	mem[2590] = 4'b1000;
	mem[2591] = 4'b1000;
	mem[2592] = 4'b1000;
	mem[2593] = 4'b1000;
	mem[2594] = 4'b0111;
	mem[2595] = 4'b1000;
	mem[2596] = 4'b0111;
	mem[2597] = 4'b0111;
	mem[2598] = 4'b1000;
	mem[2599] = 4'b1000;
	mem[2600] = 4'b0111;
	mem[2601] = 4'b1000;
	mem[2602] = 4'b1000;
	mem[2603] = 4'b1000;
	mem[2604] = 4'b1000;
	mem[2605] = 4'b0111;
	mem[2606] = 4'b0111;
	mem[2607] = 4'b0111;
	mem[2608] = 4'b0111;
	mem[2609] = 4'b0111;
	mem[2610] = 4'b0110;
	mem[2611] = 4'b0110;
	mem[2612] = 4'b0101;
	mem[2613] = 4'b0101;
	mem[2614] = 4'b0100;
	mem[2615] = 4'b0100;
	mem[2616] = 4'b0011;
	mem[2617] = 4'b0011;
	mem[2618] = 4'b0011;
	mem[2619] = 4'b0011;
	mem[2620] = 4'b0010;
	mem[2621] = 4'b0010;
	mem[2622] = 4'b0010;
	mem[2623] = 4'b0010;
	mem[2624] = 4'b0010;
	mem[2625] = 4'b0001;
	mem[2626] = 4'b0001;
	mem[2627] = 4'b0001;
	mem[2628] = 4'b0001;
	mem[2629] = 4'b0001;
	mem[2630] = 4'b0001;
	mem[2631] = 4'b0010;
	mem[2632] = 4'b0010;
	mem[2633] = 4'b0010;
	mem[2634] = 4'b0010;
	mem[2635] = 4'b1010;
	mem[2636] = 4'b1111;
	mem[2637] = 4'b1111;
	mem[2638] = 4'b1111;
	mem[2639] = 4'b1110;
	mem[2640] = 4'b1110;
	mem[2641] = 4'b1110;
	mem[2642] = 4'b1101;
	mem[2643] = 4'b1101;
	mem[2644] = 4'b1101;
	mem[2645] = 4'b1100;
	mem[2646] = 4'b1100;
	mem[2647] = 4'b1100;
	mem[2648] = 4'b1010;
	mem[2649] = 4'b1001;
	mem[2650] = 4'b1001;
	mem[2651] = 4'b1001;
	mem[2652] = 4'b1001;
	mem[2653] = 4'b1000;
	mem[2654] = 4'b0111;
	mem[2655] = 4'b0111;
	mem[2656] = 4'b0111;
	mem[2657] = 4'b0110;
	mem[2658] = 4'b0110;
	mem[2659] = 4'b0111;
	mem[2660] = 4'b0111;
	mem[2661] = 4'b0110;
	mem[2662] = 4'b0101;
	mem[2663] = 4'b0101;
	mem[2664] = 4'b0101;
	mem[2665] = 4'b0110;
	mem[2666] = 4'b0110;
	mem[2667] = 4'b0110;
	mem[2668] = 4'b0101;
	mem[2669] = 4'b0101;
	mem[2670] = 4'b0101;
	mem[2671] = 4'b0101;
	mem[2672] = 4'b0100;
	mem[2673] = 4'b0100;
	mem[2674] = 4'b0100;
	mem[2675] = 4'b0100;
	mem[2676] = 4'b0011;
	mem[2677] = 4'b0011;
	mem[2678] = 4'b0011;
	mem[2679] = 4'b0011;
	mem[2680] = 4'b0011;
	mem[2681] = 4'b0010;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b1001;
	mem[2692] = 4'b1111;
	mem[2693] = 4'b1111;
	mem[2694] = 4'b1111;
	mem[2695] = 4'b1111;
	mem[2696] = 4'b1110;
	mem[2697] = 4'b1110;
	mem[2698] = 4'b1110;
	mem[2699] = 4'b1110;
	mem[2700] = 4'b1101;
	mem[2701] = 4'b1101;
	mem[2702] = 4'b1101;
	mem[2703] = 4'b1101;
	mem[2704] = 4'b1101;
	mem[2705] = 4'b1100;
	mem[2706] = 4'b1100;
	mem[2707] = 4'b1100;
	mem[2708] = 4'b1100;
	mem[2709] = 4'b1011;
	mem[2710] = 4'b1011;
	mem[2711] = 4'b1011;
	mem[2712] = 4'b1011;
	mem[2713] = 4'b1011;
	mem[2714] = 4'b1010;
	mem[2715] = 4'b1010;
	mem[2716] = 4'b1010;
	mem[2717] = 4'b1010;
	mem[2718] = 4'b1001;
	mem[2719] = 4'b1001;
	mem[2720] = 4'b1001;
	mem[2721] = 4'b1001;
	mem[2722] = 4'b1001;
	mem[2723] = 4'b1000;
	mem[2724] = 4'b1000;
	mem[2725] = 4'b0111;
	mem[2726] = 4'b0111;
	mem[2727] = 4'b0111;
	mem[2728] = 4'b0111;
	mem[2729] = 4'b0110;
	mem[2730] = 4'b0111;
	mem[2731] = 4'b0111;
	mem[2732] = 4'b0110;
	mem[2733] = 4'b0110;
	mem[2734] = 4'b0110;
	mem[2735] = 4'b0110;
	mem[2736] = 4'b0101;
	mem[2737] = 4'b0101;
	mem[2738] = 4'b0101;
	mem[2739] = 4'b0100;
	mem[2740] = 4'b0100;
	mem[2741] = 4'b0100;
	mem[2742] = 4'b0100;
	mem[2743] = 4'b0101;
	mem[2744] = 4'b0100;
	mem[2745] = 4'b0100;
	mem[2746] = 4'b0011;
	mem[2747] = 4'b0011;
	mem[2748] = 4'b0011;
	mem[2749] = 4'b0011;
	mem[2750] = 4'b0010;
	mem[2751] = 4'b0010;
	mem[2752] = 4'b0010;
	mem[2753] = 4'b0010;
	mem[2754] = 4'b0010;
	mem[2755] = 4'b0001;
	mem[2756] = 4'b0001;
	mem[2757] = 4'b0001;
	mem[2758] = 4'b0001;
	mem[2759] = 4'b0000;
	mem[2760] = 4'b0000;
	mem[2761] = 4'b0000;
	mem[2762] = 4'b0000;
	mem[2763] = 4'b1001;
	mem[2764] = 4'b1111;
	mem[2765] = 4'b1111;
	mem[2766] = 4'b1110;
	mem[2767] = 4'b1110;
	mem[2768] = 4'b1110;
	mem[2769] = 4'b1101;
	mem[2770] = 4'b1101;
	mem[2771] = 4'b1101;
	mem[2772] = 4'b1100;
	mem[2773] = 4'b1100;
	mem[2774] = 4'b1100;
	mem[2775] = 4'b1011;
	mem[2776] = 4'b1011;
	mem[2777] = 4'b1011;
	mem[2778] = 4'b1010;
	mem[2779] = 4'b1001;
	mem[2780] = 4'b1010;
	mem[2781] = 4'b1001;
	mem[2782] = 4'b1001;
	mem[2783] = 4'b1000;
	mem[2784] = 4'b0111;
	mem[2785] = 4'b0111;
	mem[2786] = 4'b1000;
	mem[2787] = 4'b1000;
	mem[2788] = 4'b0111;
	mem[2789] = 4'b0111;
	mem[2790] = 4'b0110;
	mem[2791] = 4'b0110;
	mem[2792] = 4'b0110;
	mem[2793] = 4'b0101;
	mem[2794] = 4'b0101;
	mem[2795] = 4'b0101;
	mem[2796] = 4'b0100;
	mem[2797] = 4'b0100;
	mem[2798] = 4'b0100;
	mem[2799] = 4'b0100;
	mem[2800] = 4'b0011;
	mem[2801] = 4'b0011;
	mem[2802] = 4'b0011;
	mem[2803] = 4'b0011;
	mem[2804] = 4'b0010;
	mem[2805] = 4'b0010;
	mem[2806] = 4'b0010;
	mem[2807] = 4'b0010;
	mem[2808] = 4'b0010;
	mem[2809] = 4'b0001;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b1001;
	mem[2820] = 4'b1111;
	mem[2821] = 4'b1111;
	mem[2822] = 4'b1111;
	mem[2823] = 4'b1111;
	mem[2824] = 4'b1110;
	mem[2825] = 4'b1110;
	mem[2826] = 4'b1110;
	mem[2827] = 4'b1110;
	mem[2828] = 4'b1101;
	mem[2829] = 4'b1101;
	mem[2830] = 4'b1101;
	mem[2831] = 4'b1101;
	mem[2832] = 4'b1101;
	mem[2833] = 4'b1100;
	mem[2834] = 4'b1100;
	mem[2835] = 4'b1100;
	mem[2836] = 4'b1100;
	mem[2837] = 4'b1011;
	mem[2838] = 4'b1011;
	mem[2839] = 4'b1011;
	mem[2840] = 4'b1011;
	mem[2841] = 4'b1011;
	mem[2842] = 4'b1010;
	mem[2843] = 4'b1010;
	mem[2844] = 4'b1010;
	mem[2845] = 4'b1010;
	mem[2846] = 4'b1001;
	mem[2847] = 4'b1001;
	mem[2848] = 4'b1001;
	mem[2849] = 4'b1001;
	mem[2850] = 4'b1001;
	mem[2851] = 4'b1000;
	mem[2852] = 4'b1000;
	mem[2853] = 4'b1000;
	mem[2854] = 4'b0111;
	mem[2855] = 4'b0111;
	mem[2856] = 4'b0111;
	mem[2857] = 4'b0110;
	mem[2858] = 4'b0110;
	mem[2859] = 4'b0111;
	mem[2860] = 4'b0111;
	mem[2861] = 4'b0110;
	mem[2862] = 4'b0110;
	mem[2863] = 4'b0110;
	mem[2864] = 4'b0101;
	mem[2865] = 4'b0101;
	mem[2866] = 4'b0101;
	mem[2867] = 4'b0101;
	mem[2868] = 4'b0100;
	mem[2869] = 4'b0100;
	mem[2870] = 4'b0101;
	mem[2871] = 4'b0100;
	mem[2872] = 4'b0100;
	mem[2873] = 4'b0100;
	mem[2874] = 4'b0011;
	mem[2875] = 4'b0011;
	mem[2876] = 4'b0011;
	mem[2877] = 4'b0011;
	mem[2878] = 4'b0010;
	mem[2879] = 4'b0010;
	mem[2880] = 4'b0010;
	mem[2881] = 4'b0010;
	mem[2882] = 4'b0010;
	mem[2883] = 4'b0001;
	mem[2884] = 4'b0001;
	mem[2885] = 4'b0001;
	mem[2886] = 4'b0001;
	mem[2887] = 4'b0000;
	mem[2888] = 4'b0000;
	mem[2889] = 4'b0000;
	mem[2890] = 4'b0000;
	mem[2891] = 4'b1001;
	mem[2892] = 4'b1111;
	mem[2893] = 4'b1111;
	mem[2894] = 4'b1110;
	mem[2895] = 4'b1110;
	mem[2896] = 4'b1110;
	mem[2897] = 4'b1101;
	mem[2898] = 4'b1101;
	mem[2899] = 4'b1101;
	mem[2900] = 4'b1100;
	mem[2901] = 4'b1100;
	mem[2902] = 4'b1100;
	mem[2903] = 4'b1011;
	mem[2904] = 4'b1011;
	mem[2905] = 4'b1010;
	mem[2906] = 4'b1001;
	mem[2907] = 4'b1001;
	mem[2908] = 4'b1001;
	mem[2909] = 4'b1010;
	mem[2910] = 4'b1001;
	mem[2911] = 4'b1000;
	mem[2912] = 4'b0111;
	mem[2913] = 4'b1000;
	mem[2914] = 4'b1000;
	mem[2915] = 4'b0111;
	mem[2916] = 4'b0111;
	mem[2917] = 4'b0111;
	mem[2918] = 4'b0110;
	mem[2919] = 4'b0110;
	mem[2920] = 4'b0110;
	mem[2921] = 4'b0101;
	mem[2922] = 4'b0101;
	mem[2923] = 4'b0101;
	mem[2924] = 4'b0101;
	mem[2925] = 4'b0100;
	mem[2926] = 4'b0100;
	mem[2927] = 4'b0100;
	mem[2928] = 4'b0100;
	mem[2929] = 4'b0011;
	mem[2930] = 4'b0011;
	mem[2931] = 4'b0011;
	mem[2932] = 4'b0011;
	mem[2933] = 4'b0010;
	mem[2934] = 4'b0010;
	mem[2935] = 4'b0010;
	mem[2936] = 4'b0010;
	mem[2937] = 4'b0010;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b1001;
	mem[2948] = 4'b1111;
	mem[2949] = 4'b1111;
	mem[2950] = 4'b1111;
	mem[2951] = 4'b1111;
	mem[2952] = 4'b1110;
	mem[2953] = 4'b1110;
	mem[2954] = 4'b1110;
	mem[2955] = 4'b1110;
	mem[2956] = 4'b1101;
	mem[2957] = 4'b1101;
	mem[2958] = 4'b1101;
	mem[2959] = 4'b1101;
	mem[2960] = 4'b1101;
	mem[2961] = 4'b1100;
	mem[2962] = 4'b1100;
	mem[2963] = 4'b1100;
	mem[2964] = 4'b1100;
	mem[2965] = 4'b1011;
	mem[2966] = 4'b1011;
	mem[2967] = 4'b1011;
	mem[2968] = 4'b1011;
	mem[2969] = 4'b1011;
	mem[2970] = 4'b1010;
	mem[2971] = 4'b1010;
	mem[2972] = 4'b1010;
	mem[2973] = 4'b1010;
	mem[2974] = 4'b1001;
	mem[2975] = 4'b1001;
	mem[2976] = 4'b1001;
	mem[2977] = 4'b1001;
	mem[2978] = 4'b1001;
	mem[2979] = 4'b1000;
	mem[2980] = 4'b1000;
	mem[2981] = 4'b1000;
	mem[2982] = 4'b1000;
	mem[2983] = 4'b0111;
	mem[2984] = 4'b0110;
	mem[2985] = 4'b0110;
	mem[2986] = 4'b0110;
	mem[2987] = 4'b0110;
	mem[2988] = 4'b0111;
	mem[2989] = 4'b0110;
	mem[2990] = 4'b0110;
	mem[2991] = 4'b0110;
	mem[2992] = 4'b0101;
	mem[2993] = 4'b0101;
	mem[2994] = 4'b0101;
	mem[2995] = 4'b0101;
	mem[2996] = 4'b0101;
	mem[2997] = 4'b0101;
	mem[2998] = 4'b0101;
	mem[2999] = 4'b0100;
	mem[3000] = 4'b0100;
	mem[3001] = 4'b0100;
	mem[3002] = 4'b0011;
	mem[3003] = 4'b0011;
	mem[3004] = 4'b0011;
	mem[3005] = 4'b0011;
	mem[3006] = 4'b0010;
	mem[3007] = 4'b0010;
	mem[3008] = 4'b0010;
	mem[3009] = 4'b0010;
	mem[3010] = 4'b0010;
	mem[3011] = 4'b0001;
	mem[3012] = 4'b0001;
	mem[3013] = 4'b0001;
	mem[3014] = 4'b0001;
	mem[3015] = 4'b0000;
	mem[3016] = 4'b0000;
	mem[3017] = 4'b0000;
	mem[3018] = 4'b0000;
	mem[3019] = 4'b1001;
	mem[3020] = 4'b1111;
	mem[3021] = 4'b1111;
	mem[3022] = 4'b1110;
	mem[3023] = 4'b1110;
	mem[3024] = 4'b1110;
	mem[3025] = 4'b1101;
	mem[3026] = 4'b1101;
	mem[3027] = 4'b1101;
	mem[3028] = 4'b1100;
	mem[3029] = 4'b1100;
	mem[3030] = 4'b1100;
	mem[3031] = 4'b1011;
	mem[3032] = 4'b1010;
	mem[3033] = 4'b1001;
	mem[3034] = 4'b1001;
	mem[3035] = 4'b1001;
	mem[3036] = 4'b1010;
	mem[3037] = 4'b1010;
	mem[3038] = 4'b1001;
	mem[3039] = 4'b1001;
	mem[3040] = 4'b1001;
	mem[3041] = 4'b1001;
	mem[3042] = 4'b1000;
	mem[3043] = 4'b0111;
	mem[3044] = 4'b0111;
	mem[3045] = 4'b0111;
	mem[3046] = 4'b0110;
	mem[3047] = 4'b0110;
	mem[3048] = 4'b0110;
	mem[3049] = 4'b0110;
	mem[3050] = 4'b0101;
	mem[3051] = 4'b0101;
	mem[3052] = 4'b0101;
	mem[3053] = 4'b0101;
	mem[3054] = 4'b0100;
	mem[3055] = 4'b0100;
	mem[3056] = 4'b0100;
	mem[3057] = 4'b0100;
	mem[3058] = 4'b0011;
	mem[3059] = 4'b0011;
	mem[3060] = 4'b0011;
	mem[3061] = 4'b0011;
	mem[3062] = 4'b0011;
	mem[3063] = 4'b0010;
	mem[3064] = 4'b0010;
	mem[3065] = 4'b0010;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b1001;
	mem[3076] = 4'b1111;
	mem[3077] = 4'b1111;
	mem[3078] = 4'b1111;
	mem[3079] = 4'b1111;
	mem[3080] = 4'b1110;
	mem[3081] = 4'b1110;
	mem[3082] = 4'b1110;
	mem[3083] = 4'b1110;
	mem[3084] = 4'b1101;
	mem[3085] = 4'b1101;
	mem[3086] = 4'b1101;
	mem[3087] = 4'b1101;
	mem[3088] = 4'b1101;
	mem[3089] = 4'b1100;
	mem[3090] = 4'b1100;
	mem[3091] = 4'b1100;
	mem[3092] = 4'b1100;
	mem[3093] = 4'b1011;
	mem[3094] = 4'b1011;
	mem[3095] = 4'b1011;
	mem[3096] = 4'b1011;
	mem[3097] = 4'b1011;
	mem[3098] = 4'b1010;
	mem[3099] = 4'b1010;
	mem[3100] = 4'b1010;
	mem[3101] = 4'b1010;
	mem[3102] = 4'b1001;
	mem[3103] = 4'b1001;
	mem[3104] = 4'b1001;
	mem[3105] = 4'b1001;
	mem[3106] = 4'b1001;
	mem[3107] = 4'b1000;
	mem[3108] = 4'b1000;
	mem[3109] = 4'b1000;
	mem[3110] = 4'b1000;
	mem[3111] = 4'b1000;
	mem[3112] = 4'b0111;
	mem[3113] = 4'b0110;
	mem[3114] = 4'b0110;
	mem[3115] = 4'b0110;
	mem[3116] = 4'b0110;
	mem[3117] = 4'b0110;
	mem[3118] = 4'b0110;
	mem[3119] = 4'b0110;
	mem[3120] = 4'b0101;
	mem[3121] = 4'b0101;
	mem[3122] = 4'b0101;
	mem[3123] = 4'b0101;
	mem[3124] = 4'b0101;
	mem[3125] = 4'b0101;
	mem[3126] = 4'b0100;
	mem[3127] = 4'b0100;
	mem[3128] = 4'b0100;
	mem[3129] = 4'b0100;
	mem[3130] = 4'b0011;
	mem[3131] = 4'b0011;
	mem[3132] = 4'b0011;
	mem[3133] = 4'b0011;
	mem[3134] = 4'b0010;
	mem[3135] = 4'b0010;
	mem[3136] = 4'b0010;
	mem[3137] = 4'b0010;
	mem[3138] = 4'b0010;
	mem[3139] = 4'b0001;
	mem[3140] = 4'b0001;
	mem[3141] = 4'b0001;
	mem[3142] = 4'b0001;
	mem[3143] = 4'b0000;
	mem[3144] = 4'b0000;
	mem[3145] = 4'b0000;
	mem[3146] = 4'b0000;
	mem[3147] = 4'b1001;
	mem[3148] = 4'b1111;
	mem[3149] = 4'b1111;
	mem[3150] = 4'b1110;
	mem[3151] = 4'b1110;
	mem[3152] = 4'b1110;
	mem[3153] = 4'b1101;
	mem[3154] = 4'b1101;
	mem[3155] = 4'b1100;
	mem[3156] = 4'b1011;
	mem[3157] = 4'b1011;
	mem[3158] = 4'b1100;
	mem[3159] = 4'b1011;
	mem[3160] = 4'b1011;
	mem[3161] = 4'b1001;
	mem[3162] = 4'b1001;
	mem[3163] = 4'b1011;
	mem[3164] = 4'b1010;
	mem[3165] = 4'b1001;
	mem[3166] = 4'b1001;
	mem[3167] = 4'b1001;
	mem[3168] = 4'b1000;
	mem[3169] = 4'b1000;
	mem[3170] = 4'b1000;
	mem[3171] = 4'b0111;
	mem[3172] = 4'b0111;
	mem[3173] = 4'b0111;
	mem[3174] = 4'b0110;
	mem[3175] = 4'b0110;
	mem[3176] = 4'b0110;
	mem[3177] = 4'b0110;
	mem[3178] = 4'b0101;
	mem[3179] = 4'b0101;
	mem[3180] = 4'b0101;
	mem[3181] = 4'b0101;
	mem[3182] = 4'b0100;
	mem[3183] = 4'b0100;
	mem[3184] = 4'b0100;
	mem[3185] = 4'b0100;
	mem[3186] = 4'b0100;
	mem[3187] = 4'b0011;
	mem[3188] = 4'b0011;
	mem[3189] = 4'b0011;
	mem[3190] = 4'b0011;
	mem[3191] = 4'b0011;
	mem[3192] = 4'b0010;
	mem[3193] = 4'b0010;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b1001;
	mem[3204] = 4'b1111;
	mem[3205] = 4'b1111;
	mem[3206] = 4'b1111;
	mem[3207] = 4'b1111;
	mem[3208] = 4'b1110;
	mem[3209] = 4'b1110;
	mem[3210] = 4'b1110;
	mem[3211] = 4'b1110;
	mem[3212] = 4'b1101;
	mem[3213] = 4'b1101;
	mem[3214] = 4'b1101;
	mem[3215] = 4'b1101;
	mem[3216] = 4'b1101;
	mem[3217] = 4'b1100;
	mem[3218] = 4'b1100;
	mem[3219] = 4'b1100;
	mem[3220] = 4'b1100;
	mem[3221] = 4'b1011;
	mem[3222] = 4'b1011;
	mem[3223] = 4'b1011;
	mem[3224] = 4'b1011;
	mem[3225] = 4'b1011;
	mem[3226] = 4'b1010;
	mem[3227] = 4'b1010;
	mem[3228] = 4'b1010;
	mem[3229] = 4'b1001;
	mem[3230] = 4'b1001;
	mem[3231] = 4'b1000;
	mem[3232] = 4'b1000;
	mem[3233] = 4'b1000;
	mem[3234] = 4'b1000;
	mem[3235] = 4'b1000;
	mem[3236] = 4'b1000;
	mem[3237] = 4'b1000;
	mem[3238] = 4'b1000;
	mem[3239] = 4'b0111;
	mem[3240] = 4'b1000;
	mem[3241] = 4'b0110;
	mem[3242] = 4'b0110;
	mem[3243] = 4'b0110;
	mem[3244] = 4'b0110;
	mem[3245] = 4'b0101;
	mem[3246] = 4'b0110;
	mem[3247] = 4'b0110;
	mem[3248] = 4'b0101;
	mem[3249] = 4'b0101;
	mem[3250] = 4'b0101;
	mem[3251] = 4'b0101;
	mem[3252] = 4'b0101;
	mem[3253] = 4'b0100;
	mem[3254] = 4'b0100;
	mem[3255] = 4'b0100;
	mem[3256] = 4'b0100;
	mem[3257] = 4'b0100;
	mem[3258] = 4'b0011;
	mem[3259] = 4'b0011;
	mem[3260] = 4'b0011;
	mem[3261] = 4'b0011;
	mem[3262] = 4'b0010;
	mem[3263] = 4'b0010;
	mem[3264] = 4'b0010;
	mem[3265] = 4'b0010;
	mem[3266] = 4'b0010;
	mem[3267] = 4'b0001;
	mem[3268] = 4'b0001;
	mem[3269] = 4'b0001;
	mem[3270] = 4'b0001;
	mem[3271] = 4'b0000;
	mem[3272] = 4'b0000;
	mem[3273] = 4'b0000;
	mem[3274] = 4'b0000;
	mem[3275] = 4'b1001;
	mem[3276] = 4'b1111;
	mem[3277] = 4'b1111;
	mem[3278] = 4'b1110;
	mem[3279] = 4'b1110;
	mem[3280] = 4'b1110;
	mem[3281] = 4'b1101;
	mem[3282] = 4'b1100;
	mem[3283] = 4'b1011;
	mem[3284] = 4'b1011;
	mem[3285] = 4'b1100;
	mem[3286] = 4'b1100;
	mem[3287] = 4'b1011;
	mem[3288] = 4'b1011;
	mem[3289] = 4'b1011;
	mem[3290] = 4'b1011;
	mem[3291] = 4'b1010;
	mem[3292] = 4'b1010;
	mem[3293] = 4'b1001;
	mem[3294] = 4'b1001;
	mem[3295] = 4'b1001;
	mem[3296] = 4'b1000;
	mem[3297] = 4'b1000;
	mem[3298] = 4'b1000;
	mem[3299] = 4'b0111;
	mem[3300] = 4'b0111;
	mem[3301] = 4'b0111;
	mem[3302] = 4'b0111;
	mem[3303] = 4'b0110;
	mem[3304] = 4'b0110;
	mem[3305] = 4'b0110;
	mem[3306] = 4'b0110;
	mem[3307] = 4'b0101;
	mem[3308] = 4'b0101;
	mem[3309] = 4'b0101;
	mem[3310] = 4'b0101;
	mem[3311] = 4'b0100;
	mem[3312] = 4'b0100;
	mem[3313] = 4'b0100;
	mem[3314] = 4'b0100;
	mem[3315] = 4'b0100;
	mem[3316] = 4'b0011;
	mem[3317] = 4'b0011;
	mem[3318] = 4'b0011;
	mem[3319] = 4'b0011;
	mem[3320] = 4'b0011;
	mem[3321] = 4'b0010;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b1001;
	mem[3332] = 4'b1111;
	mem[3333] = 4'b1111;
	mem[3334] = 4'b1111;
	mem[3335] = 4'b1111;
	mem[3336] = 4'b1110;
	mem[3337] = 4'b1110;
	mem[3338] = 4'b1110;
	mem[3339] = 4'b1110;
	mem[3340] = 4'b1101;
	mem[3341] = 4'b1101;
	mem[3342] = 4'b1101;
	mem[3343] = 4'b1101;
	mem[3344] = 4'b1101;
	mem[3345] = 4'b1100;
	mem[3346] = 4'b1100;
	mem[3347] = 4'b1100;
	mem[3348] = 4'b1100;
	mem[3349] = 4'b1011;
	mem[3350] = 4'b1011;
	mem[3351] = 4'b1011;
	mem[3352] = 4'b1011;
	mem[3353] = 4'b1011;
	mem[3354] = 4'b1010;
	mem[3355] = 4'b1010;
	mem[3356] = 4'b1001;
	mem[3357] = 4'b1001;
	mem[3358] = 4'b1000;
	mem[3359] = 4'b1000;
	mem[3360] = 4'b1000;
	mem[3361] = 4'b1000;
	mem[3362] = 4'b1000;
	mem[3363] = 4'b0111;
	mem[3364] = 4'b0111;
	mem[3365] = 4'b1000;
	mem[3366] = 4'b1000;
	mem[3367] = 4'b0111;
	mem[3368] = 4'b0111;
	mem[3369] = 4'b0111;
	mem[3370] = 4'b0110;
	mem[3371] = 4'b0110;
	mem[3372] = 4'b0110;
	mem[3373] = 4'b0110;
	mem[3374] = 4'b0101;
	mem[3375] = 4'b0110;
	mem[3376] = 4'b0110;
	mem[3377] = 4'b0101;
	mem[3378] = 4'b0101;
	mem[3379] = 4'b0101;
	mem[3380] = 4'b0101;
	mem[3381] = 4'b0100;
	mem[3382] = 4'b0100;
	mem[3383] = 4'b0100;
	mem[3384] = 4'b0100;
	mem[3385] = 4'b0100;
	mem[3386] = 4'b0011;
	mem[3387] = 4'b0011;
	mem[3388] = 4'b0011;
	mem[3389] = 4'b0011;
	mem[3390] = 4'b0010;
	mem[3391] = 4'b0010;
	mem[3392] = 4'b0010;
	mem[3393] = 4'b0010;
	mem[3394] = 4'b0010;
	mem[3395] = 4'b0001;
	mem[3396] = 4'b0001;
	mem[3397] = 4'b0001;
	mem[3398] = 4'b0001;
	mem[3399] = 4'b0000;
	mem[3400] = 4'b0000;
	mem[3401] = 4'b0000;
	mem[3402] = 4'b0000;
	mem[3403] = 4'b1001;
	mem[3404] = 4'b1111;
	mem[3405] = 4'b1111;
	mem[3406] = 4'b1110;
	mem[3407] = 4'b1110;
	mem[3408] = 4'b1110;
	mem[3409] = 4'b1100;
	mem[3410] = 4'b1011;
	mem[3411] = 4'b1100;
	mem[3412] = 4'b1100;
	mem[3413] = 4'b1100;
	mem[3414] = 4'b1011;
	mem[3415] = 4'b1010;
	mem[3416] = 4'b1011;
	mem[3417] = 4'b1011;
	mem[3418] = 4'b1010;
	mem[3419] = 4'b1010;
	mem[3420] = 4'b1010;
	mem[3421] = 4'b1001;
	mem[3422] = 4'b1001;
	mem[3423] = 4'b1001;
	mem[3424] = 4'b1000;
	mem[3425] = 4'b1000;
	mem[3426] = 4'b1000;
	mem[3427] = 4'b1000;
	mem[3428] = 4'b0111;
	mem[3429] = 4'b0111;
	mem[3430] = 4'b0111;
	mem[3431] = 4'b0111;
	mem[3432] = 4'b0110;
	mem[3433] = 4'b0110;
	mem[3434] = 4'b0110;
	mem[3435] = 4'b0110;
	mem[3436] = 4'b0101;
	mem[3437] = 4'b0101;
	mem[3438] = 4'b0101;
	mem[3439] = 4'b0101;
	mem[3440] = 4'b0100;
	mem[3441] = 4'b0100;
	mem[3442] = 4'b0100;
	mem[3443] = 4'b0100;
	mem[3444] = 4'b0100;
	mem[3445] = 4'b0011;
	mem[3446] = 4'b0011;
	mem[3447] = 4'b0011;
	mem[3448] = 4'b0011;
	mem[3449] = 4'b0011;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b1001;
	mem[3460] = 4'b1111;
	mem[3461] = 4'b1111;
	mem[3462] = 4'b1111;
	mem[3463] = 4'b1111;
	mem[3464] = 4'b1110;
	mem[3465] = 4'b1110;
	mem[3466] = 4'b1110;
	mem[3467] = 4'b1110;
	mem[3468] = 4'b1101;
	mem[3469] = 4'b1101;
	mem[3470] = 4'b1101;
	mem[3471] = 4'b1101;
	mem[3472] = 4'b1101;
	mem[3473] = 4'b1100;
	mem[3474] = 4'b1100;
	mem[3475] = 4'b1100;
	mem[3476] = 4'b1100;
	mem[3477] = 4'b1011;
	mem[3478] = 4'b1011;
	mem[3479] = 4'b1011;
	mem[3480] = 4'b1011;
	mem[3481] = 4'b1011;
	mem[3482] = 4'b1010;
	mem[3483] = 4'b1001;
	mem[3484] = 4'b1001;
	mem[3485] = 4'b1001;
	mem[3486] = 4'b1000;
	mem[3487] = 4'b1000;
	mem[3488] = 4'b1000;
	mem[3489] = 4'b1000;
	mem[3490] = 4'b1000;
	mem[3491] = 4'b0111;
	mem[3492] = 4'b0111;
	mem[3493] = 4'b0111;
	mem[3494] = 4'b1000;
	mem[3495] = 4'b1000;
	mem[3496] = 4'b0111;
	mem[3497] = 4'b0111;
	mem[3498] = 4'b0111;
	mem[3499] = 4'b0110;
	mem[3500] = 4'b0110;
	mem[3501] = 4'b0110;
	mem[3502] = 4'b0101;
	mem[3503] = 4'b0101;
	mem[3504] = 4'b0110;
	mem[3505] = 4'b0101;
	mem[3506] = 4'b0101;
	mem[3507] = 4'b0101;
	mem[3508] = 4'b0101;
	mem[3509] = 4'b0100;
	mem[3510] = 4'b0100;
	mem[3511] = 4'b0100;
	mem[3512] = 4'b0100;
	mem[3513] = 4'b0100;
	mem[3514] = 4'b0011;
	mem[3515] = 4'b0011;
	mem[3516] = 4'b0011;
	mem[3517] = 4'b0011;
	mem[3518] = 4'b0010;
	mem[3519] = 4'b0010;
	mem[3520] = 4'b0010;
	mem[3521] = 4'b0010;
	mem[3522] = 4'b0010;
	mem[3523] = 4'b0001;
	mem[3524] = 4'b0001;
	mem[3525] = 4'b0001;
	mem[3526] = 4'b0001;
	mem[3527] = 4'b0000;
	mem[3528] = 4'b0000;
	mem[3529] = 4'b0000;
	mem[3530] = 4'b0000;
	mem[3531] = 4'b1001;
	mem[3532] = 4'b1111;
	mem[3533] = 4'b1111;
	mem[3534] = 4'b1110;
	mem[3535] = 4'b1110;
	mem[3536] = 4'b1101;
	mem[3537] = 4'b1100;
	mem[3538] = 4'b1101;
	mem[3539] = 4'b1101;
	mem[3540] = 4'b1100;
	mem[3541] = 4'b1011;
	mem[3542] = 4'b1010;
	mem[3543] = 4'b1010;
	mem[3544] = 4'b1001;
	mem[3545] = 4'b1011;
	mem[3546] = 4'b1010;
	mem[3547] = 4'b1010;
	mem[3548] = 4'b1010;
	mem[3549] = 4'b1001;
	mem[3550] = 4'b1001;
	mem[3551] = 4'b1001;
	mem[3552] = 4'b1001;
	mem[3553] = 4'b1000;
	mem[3554] = 4'b1000;
	mem[3555] = 4'b1000;
	mem[3556] = 4'b0111;
	mem[3557] = 4'b0111;
	mem[3558] = 4'b0111;
	mem[3559] = 4'b0111;
	mem[3560] = 4'b0110;
	mem[3561] = 4'b0110;
	mem[3562] = 4'b0110;
	mem[3563] = 4'b0110;
	mem[3564] = 4'b0110;
	mem[3565] = 4'b0101;
	mem[3566] = 4'b0101;
	mem[3567] = 4'b0101;
	mem[3568] = 4'b0101;
	mem[3569] = 4'b0100;
	mem[3570] = 4'b0100;
	mem[3571] = 4'b0100;
	mem[3572] = 4'b0100;
	mem[3573] = 4'b0100;
	mem[3574] = 4'b0100;
	mem[3575] = 4'b0011;
	mem[3576] = 4'b0011;
	mem[3577] = 4'b0011;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b1001;
	mem[3588] = 4'b1111;
	mem[3589] = 4'b1111;
	mem[3590] = 4'b1111;
	mem[3591] = 4'b1111;
	mem[3592] = 4'b1110;
	mem[3593] = 4'b1110;
	mem[3594] = 4'b1110;
	mem[3595] = 4'b1110;
	mem[3596] = 4'b1101;
	mem[3597] = 4'b1101;
	mem[3598] = 4'b1101;
	mem[3599] = 4'b1101;
	mem[3600] = 4'b1101;
	mem[3601] = 4'b1100;
	mem[3602] = 4'b1100;
	mem[3603] = 4'b1100;
	mem[3604] = 4'b1100;
	mem[3605] = 4'b1011;
	mem[3606] = 4'b1011;
	mem[3607] = 4'b1011;
	mem[3608] = 4'b1011;
	mem[3609] = 4'b1011;
	mem[3610] = 4'b1010;
	mem[3611] = 4'b1001;
	mem[3612] = 4'b1001;
	mem[3613] = 4'b1001;
	mem[3614] = 4'b1001;
	mem[3615] = 4'b1001;
	mem[3616] = 4'b1001;
	mem[3617] = 4'b1000;
	mem[3618] = 4'b1000;
	mem[3619] = 4'b0111;
	mem[3620] = 4'b0111;
	mem[3621] = 4'b0111;
	mem[3622] = 4'b0111;
	mem[3623] = 4'b1000;
	mem[3624] = 4'b0111;
	mem[3625] = 4'b0111;
	mem[3626] = 4'b0111;
	mem[3627] = 4'b0111;
	mem[3628] = 4'b0110;
	mem[3629] = 4'b0110;
	mem[3630] = 4'b0101;
	mem[3631] = 4'b0101;
	mem[3632] = 4'b0110;
	mem[3633] = 4'b0101;
	mem[3634] = 4'b0101;
	mem[3635] = 4'b0101;
	mem[3636] = 4'b0101;
	mem[3637] = 4'b0100;
	mem[3638] = 4'b0100;
	mem[3639] = 4'b0100;
	mem[3640] = 4'b0100;
	mem[3641] = 4'b0100;
	mem[3642] = 4'b0011;
	mem[3643] = 4'b0011;
	mem[3644] = 4'b0011;
	mem[3645] = 4'b0011;
	mem[3646] = 4'b0010;
	mem[3647] = 4'b0010;
	mem[3648] = 4'b0010;
	mem[3649] = 4'b0010;
	mem[3650] = 4'b0010;
	mem[3651] = 4'b0001;
	mem[3652] = 4'b0001;
	mem[3653] = 4'b0001;
	mem[3654] = 4'b0001;
	mem[3655] = 4'b0000;
	mem[3656] = 4'b0000;
	mem[3657] = 4'b0000;
	mem[3658] = 4'b0000;
	mem[3659] = 4'b1001;
	mem[3660] = 4'b1111;
	mem[3661] = 4'b1111;
	mem[3662] = 4'b1110;
	mem[3663] = 4'b1110;
	mem[3664] = 4'b1101;
	mem[3665] = 4'b1100;
	mem[3666] = 4'b1100;
	mem[3667] = 4'b1100;
	mem[3668] = 4'b1011;
	mem[3669] = 4'b1010;
	mem[3670] = 4'b1010;
	mem[3671] = 4'b1010;
	mem[3672] = 4'b1010;
	mem[3673] = 4'b1010;
	mem[3674] = 4'b1011;
	mem[3675] = 4'b1010;
	mem[3676] = 4'b1010;
	mem[3677] = 4'b1010;
	mem[3678] = 4'b1001;
	mem[3679] = 4'b1001;
	mem[3680] = 4'b1001;
	mem[3681] = 4'b1000;
	mem[3682] = 4'b1000;
	mem[3683] = 4'b1000;
	mem[3684] = 4'b1000;
	mem[3685] = 4'b0111;
	mem[3686] = 4'b0111;
	mem[3687] = 4'b0111;
	mem[3688] = 4'b0111;
	mem[3689] = 4'b0110;
	mem[3690] = 4'b0110;
	mem[3691] = 4'b0110;
	mem[3692] = 4'b0110;
	mem[3693] = 4'b0110;
	mem[3694] = 4'b0101;
	mem[3695] = 4'b0101;
	mem[3696] = 4'b0101;
	mem[3697] = 4'b0101;
	mem[3698] = 4'b0101;
	mem[3699] = 4'b0100;
	mem[3700] = 4'b0100;
	mem[3701] = 4'b0100;
	mem[3702] = 4'b0100;
	mem[3703] = 4'b0100;
	mem[3704] = 4'b0100;
	mem[3705] = 4'b0011;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b1001;
	mem[3716] = 4'b1111;
	mem[3717] = 4'b1111;
	mem[3718] = 4'b1111;
	mem[3719] = 4'b1111;
	mem[3720] = 4'b1110;
	mem[3721] = 4'b1110;
	mem[3722] = 4'b1110;
	mem[3723] = 4'b1110;
	mem[3724] = 4'b1101;
	mem[3725] = 4'b1101;
	mem[3726] = 4'b1101;
	mem[3727] = 4'b1101;
	mem[3728] = 4'b1101;
	mem[3729] = 4'b1100;
	mem[3730] = 4'b1100;
	mem[3731] = 4'b1100;
	mem[3732] = 4'b1100;
	mem[3733] = 4'b1011;
	mem[3734] = 4'b1011;
	mem[3735] = 4'b1011;
	mem[3736] = 4'b1011;
	mem[3737] = 4'b1010;
	mem[3738] = 4'b1001;
	mem[3739] = 4'b1001;
	mem[3740] = 4'b1001;
	mem[3741] = 4'b1001;
	mem[3742] = 4'b1010;
	mem[3743] = 4'b1010;
	mem[3744] = 4'b1001;
	mem[3745] = 4'b1001;
	mem[3746] = 4'b1001;
	mem[3747] = 4'b0111;
	mem[3748] = 4'b0111;
	mem[3749] = 4'b0111;
	mem[3750] = 4'b0111;
	mem[3751] = 4'b0111;
	mem[3752] = 4'b1000;
	mem[3753] = 4'b0111;
	mem[3754] = 4'b0111;
	mem[3755] = 4'b0111;
	mem[3756] = 4'b0111;
	mem[3757] = 4'b0110;
	mem[3758] = 4'b0110;
	mem[3759] = 4'b0111;
	mem[3760] = 4'b0110;
	mem[3761] = 4'b0101;
	mem[3762] = 4'b0101;
	mem[3763] = 4'b0101;
	mem[3764] = 4'b0101;
	mem[3765] = 4'b0100;
	mem[3766] = 4'b0100;
	mem[3767] = 4'b0100;
	mem[3768] = 4'b0100;
	mem[3769] = 4'b0100;
	mem[3770] = 4'b0011;
	mem[3771] = 4'b0011;
	mem[3772] = 4'b0011;
	mem[3773] = 4'b0011;
	mem[3774] = 4'b0010;
	mem[3775] = 4'b0010;
	mem[3776] = 4'b0010;
	mem[3777] = 4'b0010;
	mem[3778] = 4'b0010;
	mem[3779] = 4'b0001;
	mem[3780] = 4'b0001;
	mem[3781] = 4'b0001;
	mem[3782] = 4'b0001;
	mem[3783] = 4'b0000;
	mem[3784] = 4'b0000;
	mem[3785] = 4'b0000;
	mem[3786] = 4'b0000;
	mem[3787] = 4'b1001;
	mem[3788] = 4'b1111;
	mem[3789] = 4'b1111;
	mem[3790] = 4'b1110;
	mem[3791] = 4'b1110;
	mem[3792] = 4'b1110;
	mem[3793] = 4'b1011;
	mem[3794] = 4'b1011;
	mem[3795] = 4'b1011;
	mem[3796] = 4'b1011;
	mem[3797] = 4'b1011;
	mem[3798] = 4'b1100;
	mem[3799] = 4'b1100;
	mem[3800] = 4'b1010;
	mem[3801] = 4'b1010;
	mem[3802] = 4'b1011;
	mem[3803] = 4'b1010;
	mem[3804] = 4'b1010;
	mem[3805] = 4'b1010;
	mem[3806] = 4'b1001;
	mem[3807] = 4'b1001;
	mem[3808] = 4'b1001;
	mem[3809] = 4'b1001;
	mem[3810] = 4'b1000;
	mem[3811] = 4'b1000;
	mem[3812] = 4'b1000;
	mem[3813] = 4'b1000;
	mem[3814] = 4'b0111;
	mem[3815] = 4'b0111;
	mem[3816] = 4'b0111;
	mem[3817] = 4'b0111;
	mem[3818] = 4'b0110;
	mem[3819] = 4'b0110;
	mem[3820] = 4'b0110;
	mem[3821] = 4'b0110;
	mem[3822] = 4'b0110;
	mem[3823] = 4'b0101;
	mem[3824] = 4'b0101;
	mem[3825] = 4'b0101;
	mem[3826] = 4'b0101;
	mem[3827] = 4'b0101;
	mem[3828] = 4'b0100;
	mem[3829] = 4'b0100;
	mem[3830] = 4'b0100;
	mem[3831] = 4'b0100;
	mem[3832] = 4'b0100;
	mem[3833] = 4'b0011;
	mem[3834] = 4'b0000;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b1001;
	mem[3844] = 4'b1111;
	mem[3845] = 4'b1111;
	mem[3846] = 4'b1111;
	mem[3847] = 4'b1111;
	mem[3848] = 4'b1110;
	mem[3849] = 4'b1110;
	mem[3850] = 4'b1110;
	mem[3851] = 4'b1110;
	mem[3852] = 4'b1101;
	mem[3853] = 4'b1101;
	mem[3854] = 4'b1101;
	mem[3855] = 4'b1101;
	mem[3856] = 4'b1101;
	mem[3857] = 4'b1100;
	mem[3858] = 4'b1100;
	mem[3859] = 4'b1100;
	mem[3860] = 4'b1100;
	mem[3861] = 4'b1011;
	mem[3862] = 4'b1011;
	mem[3863] = 4'b1011;
	mem[3864] = 4'b1011;
	mem[3865] = 4'b1010;
	mem[3866] = 4'b1001;
	mem[3867] = 4'b1001;
	mem[3868] = 4'b1001;
	mem[3869] = 4'b1010;
	mem[3870] = 4'b1010;
	mem[3871] = 4'b1001;
	mem[3872] = 4'b1001;
	mem[3873] = 4'b1001;
	mem[3874] = 4'b1001;
	mem[3875] = 4'b1001;
	mem[3876] = 4'b0111;
	mem[3877] = 4'b0111;
	mem[3878] = 4'b0111;
	mem[3879] = 4'b0111;
	mem[3880] = 4'b0111;
	mem[3881] = 4'b0111;
	mem[3882] = 4'b0111;
	mem[3883] = 4'b0111;
	mem[3884] = 4'b0110;
	mem[3885] = 4'b0111;
	mem[3886] = 4'b0111;
	mem[3887] = 4'b0110;
	mem[3888] = 4'b0101;
	mem[3889] = 4'b0101;
	mem[3890] = 4'b0101;
	mem[3891] = 4'b0101;
	mem[3892] = 4'b0101;
	mem[3893] = 4'b0100;
	mem[3894] = 4'b0100;
	mem[3895] = 4'b0100;
	mem[3896] = 4'b0100;
	mem[3897] = 4'b0100;
	mem[3898] = 4'b0011;
	mem[3899] = 4'b0011;
	mem[3900] = 4'b0011;
	mem[3901] = 4'b0011;
	mem[3902] = 4'b0010;
	mem[3903] = 4'b0010;
	mem[3904] = 4'b0010;
	mem[3905] = 4'b0010;
	mem[3906] = 4'b0010;
	mem[3907] = 4'b0001;
	mem[3908] = 4'b0001;
	mem[3909] = 4'b0001;
	mem[3910] = 4'b0001;
	mem[3911] = 4'b0000;
	mem[3912] = 4'b0000;
	mem[3913] = 4'b0000;
	mem[3914] = 4'b0000;
	mem[3915] = 4'b1001;
	mem[3916] = 4'b1111;
	mem[3917] = 4'b1110;
	mem[3918] = 4'b1110;
	mem[3919] = 4'b1110;
	mem[3920] = 4'b1110;
	mem[3921] = 4'b1101;
	mem[3922] = 4'b1100;
	mem[3923] = 4'b1100;
	mem[3924] = 4'b1100;
	mem[3925] = 4'b1100;
	mem[3926] = 4'b1100;
	mem[3927] = 4'b1011;
	mem[3928] = 4'b1010;
	mem[3929] = 4'b1011;
	mem[3930] = 4'b1011;
	mem[3931] = 4'b1010;
	mem[3932] = 4'b1010;
	mem[3933] = 4'b1010;
	mem[3934] = 4'b1001;
	mem[3935] = 4'b1001;
	mem[3936] = 4'b1001;
	mem[3937] = 4'b1001;
	mem[3938] = 4'b1000;
	mem[3939] = 4'b1000;
	mem[3940] = 4'b1000;
	mem[3941] = 4'b1000;
	mem[3942] = 4'b0111;
	mem[3943] = 4'b0111;
	mem[3944] = 4'b0111;
	mem[3945] = 4'b0111;
	mem[3946] = 4'b0111;
	mem[3947] = 4'b0110;
	mem[3948] = 4'b0110;
	mem[3949] = 4'b0110;
	mem[3950] = 4'b0110;
	mem[3951] = 4'b0110;
	mem[3952] = 4'b0101;
	mem[3953] = 4'b0101;
	mem[3954] = 4'b0101;
	mem[3955] = 4'b0101;
	mem[3956] = 4'b0101;
	mem[3957] = 4'b0100;
	mem[3958] = 4'b0100;
	mem[3959] = 4'b0100;
	mem[3960] = 4'b0100;
	mem[3961] = 4'b0100;
	mem[3962] = 4'b0001;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b1001;
	mem[3972] = 4'b1111;
	mem[3973] = 4'b1111;
	mem[3974] = 4'b1111;
	mem[3975] = 4'b1111;
	mem[3976] = 4'b1110;
	mem[3977] = 4'b1110;
	mem[3978] = 4'b1110;
	mem[3979] = 4'b1110;
	mem[3980] = 4'b1101;
	mem[3981] = 4'b1101;
	mem[3982] = 4'b1101;
	mem[3983] = 4'b1101;
	mem[3984] = 4'b1101;
	mem[3985] = 4'b1100;
	mem[3986] = 4'b1100;
	mem[3987] = 4'b1100;
	mem[3988] = 4'b1100;
	mem[3989] = 4'b1011;
	mem[3990] = 4'b1011;
	mem[3991] = 4'b1011;
	mem[3992] = 4'b1011;
	mem[3993] = 4'b1010;
	mem[3994] = 4'b1001;
	mem[3995] = 4'b1001;
	mem[3996] = 4'b1001;
	mem[3997] = 4'b1010;
	mem[3998] = 4'b1001;
	mem[3999] = 4'b1001;
	mem[4000] = 4'b1001;
	mem[4001] = 4'b1001;
	mem[4002] = 4'b1001;
	mem[4003] = 4'b1000;
	mem[4004] = 4'b1000;
	mem[4005] = 4'b0111;
	mem[4006] = 4'b0111;
	mem[4007] = 4'b0111;
	mem[4008] = 4'b0111;
	mem[4009] = 4'b0111;
	mem[4010] = 4'b0111;
	mem[4011] = 4'b0111;
	mem[4012] = 4'b0110;
	mem[4013] = 4'b0110;
	mem[4014] = 4'b0110;
	mem[4015] = 4'b0110;
	mem[4016] = 4'b0101;
	mem[4017] = 4'b0101;
	mem[4018] = 4'b0101;
	mem[4019] = 4'b0101;
	mem[4020] = 4'b0101;
	mem[4021] = 4'b0100;
	mem[4022] = 4'b0100;
	mem[4023] = 4'b0100;
	mem[4024] = 4'b0100;
	mem[4025] = 4'b0100;
	mem[4026] = 4'b0011;
	mem[4027] = 4'b0011;
	mem[4028] = 4'b0011;
	mem[4029] = 4'b0011;
	mem[4030] = 4'b0010;
	mem[4031] = 4'b0010;
	mem[4032] = 4'b0010;
	mem[4033] = 4'b0010;
	mem[4034] = 4'b0010;
	mem[4035] = 4'b0001;
	mem[4036] = 4'b0001;
	mem[4037] = 4'b0001;
	mem[4038] = 4'b0001;
	mem[4039] = 4'b0000;
	mem[4040] = 4'b0000;
	mem[4041] = 4'b0000;
	mem[4042] = 4'b0000;
	mem[4043] = 4'b1001;
	mem[4044] = 4'b1110;
	mem[4045] = 4'b1101;
	mem[4046] = 4'b1101;
	mem[4047] = 4'b1101;
	mem[4048] = 4'b1110;
	mem[4049] = 4'b1101;
	mem[4050] = 4'b1101;
	mem[4051] = 4'b1101;
	mem[4052] = 4'b1100;
	mem[4053] = 4'b1011;
	mem[4054] = 4'b1011;
	mem[4055] = 4'b1010;
	mem[4056] = 4'b1010;
	mem[4057] = 4'b1011;
	mem[4058] = 4'b1011;
	mem[4059] = 4'b1010;
	mem[4060] = 4'b1010;
	mem[4061] = 4'b1010;
	mem[4062] = 4'b1010;
	mem[4063] = 4'b1001;
	mem[4064] = 4'b1001;
	mem[4065] = 4'b1001;
	mem[4066] = 4'b1001;
	mem[4067] = 4'b1000;
	mem[4068] = 4'b1000;
	mem[4069] = 4'b1000;
	mem[4070] = 4'b1000;
	mem[4071] = 4'b0111;
	mem[4072] = 4'b0111;
	mem[4073] = 4'b0111;
	mem[4074] = 4'b0111;
	mem[4075] = 4'b0111;
	mem[4076] = 4'b0110;
	mem[4077] = 4'b0110;
	mem[4078] = 4'b0110;
	mem[4079] = 4'b0110;
	mem[4080] = 4'b0110;
	mem[4081] = 4'b0101;
	mem[4082] = 4'b0101;
	mem[4083] = 4'b0101;
	mem[4084] = 4'b0101;
	mem[4085] = 4'b0101;
	mem[4086] = 4'b0101;
	mem[4087] = 4'b0100;
	mem[4088] = 4'b0100;
	mem[4089] = 4'b0100;
	mem[4090] = 4'b0001;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

module rom_3b (
	input clock,
	input [11:0] address,
	output reg [3:0] data_out
);

reg [3:0] mem [0:4095];

always @(posedge clock) begin
	data_out <= mem[address];
end

initial begin
	mem[0] = 4'b0000;
	mem[1] = 4'b0000;
	mem[2] = 4'b0000;
	mem[3] = 4'b0110;
	mem[4] = 4'b1001;
	mem[5] = 4'b1001;
	mem[6] = 4'b1001;
	mem[7] = 4'b1001;
	mem[8] = 4'b1001;
	mem[9] = 4'b1001;
	mem[10] = 4'b1001;
	mem[11] = 4'b1001;
	mem[12] = 4'b1001;
	mem[13] = 4'b1001;
	mem[14] = 4'b1001;
	mem[15] = 4'b1001;
	mem[16] = 4'b1001;
	mem[17] = 4'b1001;
	mem[18] = 4'b1001;
	mem[19] = 4'b1000;
	mem[20] = 4'b1001;
	mem[21] = 4'b1001;
	mem[22] = 4'b1001;
	mem[23] = 4'b1001;
	mem[24] = 4'b1000;
	mem[25] = 4'b1000;
	mem[26] = 4'b1000;
	mem[27] = 4'b1000;
	mem[28] = 4'b1000;
	mem[29] = 4'b1001;
	mem[30] = 4'b1000;
	mem[31] = 4'b1000;
	mem[32] = 4'b1000;
	mem[33] = 4'b1000;
	mem[34] = 4'b1000;
	mem[35] = 4'b1000;
	mem[36] = 4'b1000;
	mem[37] = 4'b1000;
	mem[38] = 4'b0111;
	mem[39] = 4'b0111;
	mem[40] = 4'b0111;
	mem[41] = 4'b1000;
	mem[42] = 4'b1000;
	mem[43] = 4'b1000;
	mem[44] = 4'b1000;
	mem[45] = 4'b1000;
	mem[46] = 4'b1000;
	mem[47] = 4'b1000;
	mem[48] = 4'b1000;
	mem[49] = 4'b1000;
	mem[50] = 4'b1000;
	mem[51] = 4'b1000;
	mem[52] = 4'b0111;
	mem[53] = 4'b1000;
	mem[54] = 4'b1000;
	mem[55] = 4'b1000;
	mem[56] = 4'b1000;
	mem[57] = 4'b0111;
	mem[58] = 4'b0111;
	mem[59] = 4'b0111;
	mem[60] = 4'b0111;
	mem[61] = 4'b0111;
	mem[62] = 4'b0111;
	mem[63] = 4'b0111;
	mem[64] = 4'b0111;
	mem[65] = 4'b0111;
	mem[66] = 4'b0111;
	mem[67] = 4'b0111;
	mem[68] = 4'b0111;
	mem[69] = 4'b0110;
	mem[70] = 4'b0011;
	mem[71] = 4'b0000;
	mem[72] = 4'b0000;
	mem[73] = 4'b0000;
	mem[74] = 4'b0000;
	mem[75] = 4'b0101;
	mem[76] = 4'b1000;
	mem[77] = 4'b1000;
	mem[78] = 4'b1000;
	mem[79] = 4'b1000;
	mem[80] = 4'b1000;
	mem[81] = 4'b1000;
	mem[82] = 4'b1000;
	mem[83] = 4'b1000;
	mem[84] = 4'b0111;
	mem[85] = 4'b0111;
	mem[86] = 4'b0111;
	mem[87] = 4'b1000;
	mem[88] = 4'b1000;
	mem[89] = 4'b0111;
	mem[90] = 4'b0111;
	mem[91] = 4'b0111;
	mem[92] = 4'b0111;
	mem[93] = 4'b0111;
	mem[94] = 4'b0111;
	mem[95] = 4'b0110;
	mem[96] = 4'b0110;
	mem[97] = 4'b0110;
	mem[98] = 4'b0110;
	mem[99] = 4'b0110;
	mem[100] = 4'b0110;
	mem[101] = 4'b0110;
	mem[102] = 4'b0110;
	mem[103] = 4'b0110;
	mem[104] = 4'b0101;
	mem[105] = 4'b0101;
	mem[106] = 4'b0101;
	mem[107] = 4'b0101;
	mem[108] = 4'b0101;
	mem[109] = 4'b0101;
	mem[110] = 4'b0101;
	mem[111] = 4'b0101;
	mem[112] = 4'b0101;
	mem[113] = 4'b0101;
	mem[114] = 4'b0101;
	mem[115] = 4'b0101;
	mem[116] = 4'b0101;
	mem[117] = 4'b0101;
	mem[118] = 4'b0101;
	mem[119] = 4'b0100;
	mem[120] = 4'b0100;
	mem[121] = 4'b0100;
	mem[122] = 4'b0001;
	mem[123] = 4'b0000;
	mem[124] = 4'b0000;
	mem[125] = 4'b0000;
	mem[126] = 4'b0000;
	mem[127] = 4'b0000;
	mem[128] = 4'b0000;
	mem[129] = 4'b0000;
	mem[130] = 4'b0000;
	mem[131] = 4'b0000;
	mem[132] = 4'b0000;
	mem[133] = 4'b0000;
	mem[134] = 4'b0000;
	mem[135] = 4'b0000;
	mem[136] = 4'b0000;
	mem[137] = 4'b0001;
	mem[138] = 4'b0001;
	mem[139] = 4'b0001;
	mem[140] = 4'b0001;
	mem[141] = 4'b0001;
	mem[142] = 4'b0010;
	mem[143] = 4'b0011;
	mem[144] = 4'b0011;
	mem[145] = 4'b0011;
	mem[146] = 4'b0011;
	mem[147] = 4'b0011;
	mem[148] = 4'b0100;
	mem[149] = 4'b0100;
	mem[150] = 4'b0100;
	mem[151] = 4'b0100;
	mem[152] = 4'b0100;
	mem[153] = 4'b0101;
	mem[154] = 4'b0101;
	mem[155] = 4'b0101;
	mem[156] = 4'b0110;
	mem[157] = 4'b0110;
	mem[158] = 4'b0110;
	mem[159] = 4'b0111;
	mem[160] = 4'b1000;
	mem[161] = 4'b1000;
	mem[162] = 4'b1000;
	mem[163] = 4'b1000;
	mem[164] = 4'b1000;
	mem[165] = 4'b1001;
	mem[166] = 4'b1000;
	mem[167] = 4'b1000;
	mem[168] = 4'b1000;
	mem[169] = 4'b1001;
	mem[170] = 4'b1010;
	mem[171] = 4'b1011;
	mem[172] = 4'b1011;
	mem[173] = 4'b1011;
	mem[174] = 4'b1011;
	mem[175] = 4'b1011;
	mem[176] = 4'b1100;
	mem[177] = 4'b1100;
	mem[178] = 4'b1100;
	mem[179] = 4'b1100;
	mem[180] = 4'b1100;
	mem[181] = 4'b1101;
	mem[182] = 4'b1110;
	mem[183] = 4'b1110;
	mem[184] = 4'b1110;
	mem[185] = 4'b1110;
	mem[186] = 4'b1110;
	mem[187] = 4'b1111;
	mem[188] = 4'b1111;
	mem[189] = 4'b1111;
	mem[190] = 4'b1111;
	mem[191] = 4'b1111;
	mem[192] = 4'b1111;
	mem[193] = 4'b1111;
	mem[194] = 4'b1111;
	mem[195] = 4'b1111;
	mem[196] = 4'b1111;
	mem[197] = 4'b1111;
	mem[198] = 4'b0110;
	mem[199] = 4'b0000;
	mem[200] = 4'b0000;
	mem[201] = 4'b0000;
	mem[202] = 4'b0000;
	mem[203] = 4'b0000;
	mem[204] = 4'b0001;
	mem[205] = 4'b0001;
	mem[206] = 4'b0001;
	mem[207] = 4'b0000;
	mem[208] = 4'b0000;
	mem[209] = 4'b0001;
	mem[210] = 4'b0001;
	mem[211] = 4'b0000;
	mem[212] = 4'b0001;
	mem[213] = 4'b0010;
	mem[214] = 4'b0010;
	mem[215] = 4'b0010;
	mem[216] = 4'b0001;
	mem[217] = 4'b0001;
	mem[218] = 4'b0001;
	mem[219] = 4'b0001;
	mem[220] = 4'b0001;
	mem[221] = 4'b0001;
	mem[222] = 4'b0010;
	mem[223] = 4'b0010;
	mem[224] = 4'b0010;
	mem[225] = 4'b0010;
	mem[226] = 4'b0010;
	mem[227] = 4'b0010;
	mem[228] = 4'b0010;
	mem[229] = 4'b0010;
	mem[230] = 4'b0010;
	mem[231] = 4'b0011;
	mem[232] = 4'b0011;
	mem[233] = 4'b0011;
	mem[234] = 4'b0011;
	mem[235] = 4'b0011;
	mem[236] = 4'b0011;
	mem[237] = 4'b0011;
	mem[238] = 4'b0011;
	mem[239] = 4'b0011;
	mem[240] = 4'b0100;
	mem[241] = 4'b0100;
	mem[242] = 4'b0100;
	mem[243] = 4'b0100;
	mem[244] = 4'b0100;
	mem[245] = 4'b0100;
	mem[246] = 4'b0100;
	mem[247] = 4'b0100;
	mem[248] = 4'b0100;
	mem[249] = 4'b0100;
	mem[250] = 4'b0001;
	mem[251] = 4'b0000;
	mem[252] = 4'b0000;
	mem[253] = 4'b0000;
	mem[254] = 4'b0000;
	mem[255] = 4'b0000;
	mem[256] = 4'b0000;
	mem[257] = 4'b0000;
	mem[258] = 4'b0000;
	mem[259] = 4'b0000;
	mem[260] = 4'b0000;
	mem[261] = 4'b0000;
	mem[262] = 4'b0000;
	mem[263] = 4'b0000;
	mem[264] = 4'b0000;
	mem[265] = 4'b0001;
	mem[266] = 4'b0001;
	mem[267] = 4'b0001;
	mem[268] = 4'b0001;
	mem[269] = 4'b0001;
	mem[270] = 4'b0010;
	mem[271] = 4'b0011;
	mem[272] = 4'b0011;
	mem[273] = 4'b0011;
	mem[274] = 4'b0011;
	mem[275] = 4'b0011;
	mem[276] = 4'b0100;
	mem[277] = 4'b0100;
	mem[278] = 4'b0100;
	mem[279] = 4'b0100;
	mem[280] = 4'b0100;
	mem[281] = 4'b0101;
	mem[282] = 4'b0101;
	mem[283] = 4'b0101;
	mem[284] = 4'b0101;
	mem[285] = 4'b0110;
	mem[286] = 4'b0110;
	mem[287] = 4'b0111;
	mem[288] = 4'b1000;
	mem[289] = 4'b1000;
	mem[290] = 4'b1000;
	mem[291] = 4'b1000;
	mem[292] = 4'b1000;
	mem[293] = 4'b1000;
	mem[294] = 4'b1000;
	mem[295] = 4'b1000;
	mem[296] = 4'b1001;
	mem[297] = 4'b1001;
	mem[298] = 4'b1010;
	mem[299] = 4'b1011;
	mem[300] = 4'b1011;
	mem[301] = 4'b1011;
	mem[302] = 4'b1011;
	mem[303] = 4'b1011;
	mem[304] = 4'b1100;
	mem[305] = 4'b1100;
	mem[306] = 4'b1100;
	mem[307] = 4'b1100;
	mem[308] = 4'b1100;
	mem[309] = 4'b1101;
	mem[310] = 4'b1110;
	mem[311] = 4'b1110;
	mem[312] = 4'b1110;
	mem[313] = 4'b1110;
	mem[314] = 4'b1110;
	mem[315] = 4'b1111;
	mem[316] = 4'b1111;
	mem[317] = 4'b1111;
	mem[318] = 4'b1111;
	mem[319] = 4'b1111;
	mem[320] = 4'b1111;
	mem[321] = 4'b1111;
	mem[322] = 4'b1111;
	mem[323] = 4'b1111;
	mem[324] = 4'b1111;
	mem[325] = 4'b1111;
	mem[326] = 4'b0110;
	mem[327] = 4'b0000;
	mem[328] = 4'b0000;
	mem[329] = 4'b0000;
	mem[330] = 4'b0000;
	mem[331] = 4'b0000;
	mem[332] = 4'b0001;
	mem[333] = 4'b0000;
	mem[334] = 4'b0000;
	mem[335] = 4'b0001;
	mem[336] = 4'b0001;
	mem[337] = 4'b0001;
	mem[338] = 4'b0001;
	mem[339] = 4'b0001;
	mem[340] = 4'b0001;
	mem[341] = 4'b0001;
	mem[342] = 4'b0001;
	mem[343] = 4'b0001;
	mem[344] = 4'b0001;
	mem[345] = 4'b0001;
	mem[346] = 4'b0001;
	mem[347] = 4'b0010;
	mem[348] = 4'b0010;
	mem[349] = 4'b0010;
	mem[350] = 4'b0010;
	mem[351] = 4'b0010;
	mem[352] = 4'b0010;
	mem[353] = 4'b0010;
	mem[354] = 4'b0010;
	mem[355] = 4'b0010;
	mem[356] = 4'b0011;
	mem[357] = 4'b0011;
	mem[358] = 4'b0011;
	mem[359] = 4'b0011;
	mem[360] = 4'b0011;
	mem[361] = 4'b0011;
	mem[362] = 4'b0011;
	mem[363] = 4'b0011;
	mem[364] = 4'b0011;
	mem[365] = 4'b0011;
	mem[366] = 4'b0100;
	mem[367] = 4'b0100;
	mem[368] = 4'b0100;
	mem[369] = 4'b0100;
	mem[370] = 4'b0100;
	mem[371] = 4'b0100;
	mem[372] = 4'b0100;
	mem[373] = 4'b0100;
	mem[374] = 4'b0100;
	mem[375] = 4'b0101;
	mem[376] = 4'b0101;
	mem[377] = 4'b0101;
	mem[378] = 4'b0001;
	mem[379] = 4'b0000;
	mem[380] = 4'b0000;
	mem[381] = 4'b0000;
	mem[382] = 4'b0000;
	mem[383] = 4'b0000;
	mem[384] = 4'b0000;
	mem[385] = 4'b0000;
	mem[386] = 4'b0000;
	mem[387] = 4'b0000;
	mem[388] = 4'b0000;
	mem[389] = 4'b0000;
	mem[390] = 4'b0000;
	mem[391] = 4'b0000;
	mem[392] = 4'b0000;
	mem[393] = 4'b0001;
	mem[394] = 4'b0001;
	mem[395] = 4'b0001;
	mem[396] = 4'b0001;
	mem[397] = 4'b0001;
	mem[398] = 4'b0010;
	mem[399] = 4'b0011;
	mem[400] = 4'b0011;
	mem[401] = 4'b0011;
	mem[402] = 4'b0011;
	mem[403] = 4'b0011;
	mem[404] = 4'b0100;
	mem[405] = 4'b0100;
	mem[406] = 4'b0100;
	mem[407] = 4'b0100;
	mem[408] = 4'b0100;
	mem[409] = 4'b0101;
	mem[410] = 4'b0101;
	mem[411] = 4'b0101;
	mem[412] = 4'b0101;
	mem[413] = 4'b0101;
	mem[414] = 4'b0110;
	mem[415] = 4'b0111;
	mem[416] = 4'b1000;
	mem[417] = 4'b1000;
	mem[418] = 4'b1000;
	mem[419] = 4'b1000;
	mem[420] = 4'b1000;
	mem[421] = 4'b1000;
	mem[422] = 4'b1000;
	mem[423] = 4'b1000;
	mem[424] = 4'b1001;
	mem[425] = 4'b1001;
	mem[426] = 4'b1010;
	mem[427] = 4'b1011;
	mem[428] = 4'b1011;
	mem[429] = 4'b1011;
	mem[430] = 4'b1011;
	mem[431] = 4'b1011;
	mem[432] = 4'b1100;
	mem[433] = 4'b1100;
	mem[434] = 4'b1100;
	mem[435] = 4'b1100;
	mem[436] = 4'b1100;
	mem[437] = 4'b1101;
	mem[438] = 4'b1110;
	mem[439] = 4'b1110;
	mem[440] = 4'b1110;
	mem[441] = 4'b1110;
	mem[442] = 4'b1110;
	mem[443] = 4'b1111;
	mem[444] = 4'b1111;
	mem[445] = 4'b1111;
	mem[446] = 4'b1111;
	mem[447] = 4'b1111;
	mem[448] = 4'b1111;
	mem[449] = 4'b1111;
	mem[450] = 4'b1111;
	mem[451] = 4'b1111;
	mem[452] = 4'b1111;
	mem[453] = 4'b1111;
	mem[454] = 4'b0110;
	mem[455] = 4'b0000;
	mem[456] = 4'b0000;
	mem[457] = 4'b0000;
	mem[458] = 4'b0000;
	mem[459] = 4'b0001;
	mem[460] = 4'b0001;
	mem[461] = 4'b0000;
	mem[462] = 4'b0000;
	mem[463] = 4'b0001;
	mem[464] = 4'b0001;
	mem[465] = 4'b0001;
	mem[466] = 4'b0001;
	mem[467] = 4'b0010;
	mem[468] = 4'b0001;
	mem[469] = 4'b0001;
	mem[470] = 4'b0001;
	mem[471] = 4'b0001;
	mem[472] = 4'b0001;
	mem[473] = 4'b0010;
	mem[474] = 4'b0010;
	mem[475] = 4'b0010;
	mem[476] = 4'b0010;
	mem[477] = 4'b0010;
	mem[478] = 4'b0010;
	mem[479] = 4'b0010;
	mem[480] = 4'b0010;
	mem[481] = 4'b0010;
	mem[482] = 4'b0011;
	mem[483] = 4'b0011;
	mem[484] = 4'b0011;
	mem[485] = 4'b0011;
	mem[486] = 4'b0011;
	mem[487] = 4'b0011;
	mem[488] = 4'b0011;
	mem[489] = 4'b0011;
	mem[490] = 4'b0011;
	mem[491] = 4'b0100;
	mem[492] = 4'b0100;
	mem[493] = 4'b0100;
	mem[494] = 4'b0100;
	mem[495] = 4'b0100;
	mem[496] = 4'b0100;
	mem[497] = 4'b0100;
	mem[498] = 4'b0100;
	mem[499] = 4'b0100;
	mem[500] = 4'b0101;
	mem[501] = 4'b0101;
	mem[502] = 4'b0101;
	mem[503] = 4'b0101;
	mem[504] = 4'b0101;
	mem[505] = 4'b0101;
	mem[506] = 4'b0001;
	mem[507] = 4'b0000;
	mem[508] = 4'b0000;
	mem[509] = 4'b0000;
	mem[510] = 4'b0000;
	mem[511] = 4'b0000;
	mem[512] = 4'b0000;
	mem[513] = 4'b0000;
	mem[514] = 4'b0000;
	mem[515] = 4'b0000;
	mem[516] = 4'b0000;
	mem[517] = 4'b0000;
	mem[518] = 4'b0000;
	mem[519] = 4'b0000;
	mem[520] = 4'b0000;
	mem[521] = 4'b0001;
	mem[522] = 4'b0001;
	mem[523] = 4'b0001;
	mem[524] = 4'b0001;
	mem[525] = 4'b0001;
	mem[526] = 4'b0010;
	mem[527] = 4'b0011;
	mem[528] = 4'b0011;
	mem[529] = 4'b0011;
	mem[530] = 4'b0011;
	mem[531] = 4'b0011;
	mem[532] = 4'b0100;
	mem[533] = 4'b0100;
	mem[534] = 4'b0100;
	mem[535] = 4'b0100;
	mem[536] = 4'b0100;
	mem[537] = 4'b0101;
	mem[538] = 4'b0110;
	mem[539] = 4'b0101;
	mem[540] = 4'b0101;
	mem[541] = 4'b0101;
	mem[542] = 4'b0101;
	mem[543] = 4'b0111;
	mem[544] = 4'b1000;
	mem[545] = 4'b1000;
	mem[546] = 4'b0111;
	mem[547] = 4'b0111;
	mem[548] = 4'b0111;
	mem[549] = 4'b1000;
	mem[550] = 4'b1000;
	mem[551] = 4'b1000;
	mem[552] = 4'b1010;
	mem[553] = 4'b1001;
	mem[554] = 4'b1010;
	mem[555] = 4'b1011;
	mem[556] = 4'b1011;
	mem[557] = 4'b1011;
	mem[558] = 4'b1011;
	mem[559] = 4'b1011;
	mem[560] = 4'b1100;
	mem[561] = 4'b1100;
	mem[562] = 4'b1100;
	mem[563] = 4'b1100;
	mem[564] = 4'b1100;
	mem[565] = 4'b1101;
	mem[566] = 4'b1110;
	mem[567] = 4'b1110;
	mem[568] = 4'b1110;
	mem[569] = 4'b1110;
	mem[570] = 4'b1110;
	mem[571] = 4'b1111;
	mem[572] = 4'b1111;
	mem[573] = 4'b1111;
	mem[574] = 4'b1111;
	mem[575] = 4'b1111;
	mem[576] = 4'b1111;
	mem[577] = 4'b1111;
	mem[578] = 4'b1111;
	mem[579] = 4'b1111;
	mem[580] = 4'b1111;
	mem[581] = 4'b1111;
	mem[582] = 4'b0110;
	mem[583] = 4'b0000;
	mem[584] = 4'b0000;
	mem[585] = 4'b0001;
	mem[586] = 4'b0001;
	mem[587] = 4'b0001;
	mem[588] = 4'b0001;
	mem[589] = 4'b0001;
	mem[590] = 4'b0001;
	mem[591] = 4'b0001;
	mem[592] = 4'b0001;
	mem[593] = 4'b0010;
	mem[594] = 4'b0001;
	mem[595] = 4'b0010;
	mem[596] = 4'b0010;
	mem[597] = 4'b0001;
	mem[598] = 4'b0010;
	mem[599] = 4'b0010;
	mem[600] = 4'b0010;
	mem[601] = 4'b0010;
	mem[602] = 4'b0010;
	mem[603] = 4'b0010;
	mem[604] = 4'b0010;
	mem[605] = 4'b0010;
	mem[606] = 4'b0010;
	mem[607] = 4'b0011;
	mem[608] = 4'b0011;
	mem[609] = 4'b0011;
	mem[610] = 4'b0011;
	mem[611] = 4'b0011;
	mem[612] = 4'b0011;
	mem[613] = 4'b0011;
	mem[614] = 4'b0011;
	mem[615] = 4'b0011;
	mem[616] = 4'b0100;
	mem[617] = 4'b0100;
	mem[618] = 4'b0100;
	mem[619] = 4'b0100;
	mem[620] = 4'b0100;
	mem[621] = 4'b0100;
	mem[622] = 4'b0100;
	mem[623] = 4'b0100;
	mem[624] = 4'b0100;
	mem[625] = 4'b0100;
	mem[626] = 4'b0101;
	mem[627] = 4'b0101;
	mem[628] = 4'b0101;
	mem[629] = 4'b0101;
	mem[630] = 4'b0101;
	mem[631] = 4'b0101;
	mem[632] = 4'b0101;
	mem[633] = 4'b0101;
	mem[634] = 4'b0001;
	mem[635] = 4'b0000;
	mem[636] = 4'b0000;
	mem[637] = 4'b0000;
	mem[638] = 4'b0000;
	mem[639] = 4'b0000;
	mem[640] = 4'b0000;
	mem[641] = 4'b0000;
	mem[642] = 4'b0000;
	mem[643] = 4'b0000;
	mem[644] = 4'b0000;
	mem[645] = 4'b0000;
	mem[646] = 4'b0000;
	mem[647] = 4'b0000;
	mem[648] = 4'b0000;
	mem[649] = 4'b0001;
	mem[650] = 4'b0001;
	mem[651] = 4'b0001;
	mem[652] = 4'b0001;
	mem[653] = 4'b0001;
	mem[654] = 4'b0010;
	mem[655] = 4'b0011;
	mem[656] = 4'b0011;
	mem[657] = 4'b0011;
	mem[658] = 4'b0011;
	mem[659] = 4'b0011;
	mem[660] = 4'b0100;
	mem[661] = 4'b0100;
	mem[662] = 4'b0100;
	mem[663] = 4'b0101;
	mem[664] = 4'b0100;
	mem[665] = 4'b0101;
	mem[666] = 4'b0110;
	mem[667] = 4'b0101;
	mem[668] = 4'b0101;
	mem[669] = 4'b0101;
	mem[670] = 4'b0101;
	mem[671] = 4'b0110;
	mem[672] = 4'b0111;
	mem[673] = 4'b0111;
	mem[674] = 4'b0111;
	mem[675] = 4'b0111;
	mem[676] = 4'b0111;
	mem[677] = 4'b1000;
	mem[678] = 4'b1000;
	mem[679] = 4'b1001;
	mem[680] = 4'b1001;
	mem[681] = 4'b1001;
	mem[682] = 4'b1010;
	mem[683] = 4'b1011;
	mem[684] = 4'b1011;
	mem[685] = 4'b1011;
	mem[686] = 4'b1011;
	mem[687] = 4'b1011;
	mem[688] = 4'b1100;
	mem[689] = 4'b1100;
	mem[690] = 4'b1100;
	mem[691] = 4'b1100;
	mem[692] = 4'b1100;
	mem[693] = 4'b1101;
	mem[694] = 4'b1110;
	mem[695] = 4'b1110;
	mem[696] = 4'b1110;
	mem[697] = 4'b1110;
	mem[698] = 4'b1110;
	mem[699] = 4'b1111;
	mem[700] = 4'b1111;
	mem[701] = 4'b1111;
	mem[702] = 4'b1111;
	mem[703] = 4'b1111;
	mem[704] = 4'b1111;
	mem[705] = 4'b1111;
	mem[706] = 4'b1111;
	mem[707] = 4'b1111;
	mem[708] = 4'b1111;
	mem[709] = 4'b1111;
	mem[710] = 4'b0110;
	mem[711] = 4'b0000;
	mem[712] = 4'b0000;
	mem[713] = 4'b0000;
	mem[714] = 4'b0001;
	mem[715] = 4'b0001;
	mem[716] = 4'b0001;
	mem[717] = 4'b0010;
	mem[718] = 4'b0001;
	mem[719] = 4'b0001;
	mem[720] = 4'b0001;
	mem[721] = 4'b0001;
	mem[722] = 4'b0010;
	mem[723] = 4'b0011;
	mem[724] = 4'b0010;
	mem[725] = 4'b0010;
	mem[726] = 4'b0010;
	mem[727] = 4'b0010;
	mem[728] = 4'b0010;
	mem[729] = 4'b0010;
	mem[730] = 4'b0010;
	mem[731] = 4'b0010;
	mem[732] = 4'b0010;
	mem[733] = 4'b0011;
	mem[734] = 4'b0011;
	mem[735] = 4'b0011;
	mem[736] = 4'b0011;
	mem[737] = 4'b0011;
	mem[738] = 4'b0011;
	mem[739] = 4'b0011;
	mem[740] = 4'b0011;
	mem[741] = 4'b0011;
	mem[742] = 4'b0100;
	mem[743] = 4'b0100;
	mem[744] = 4'b0100;
	mem[745] = 4'b0100;
	mem[746] = 4'b0100;
	mem[747] = 4'b0100;
	mem[748] = 4'b0100;
	mem[749] = 4'b0100;
	mem[750] = 4'b0100;
	mem[751] = 4'b0101;
	mem[752] = 4'b0101;
	mem[753] = 4'b0101;
	mem[754] = 4'b0101;
	mem[755] = 4'b0101;
	mem[756] = 4'b0101;
	mem[757] = 4'b0101;
	mem[758] = 4'b0101;
	mem[759] = 4'b0101;
	mem[760] = 4'b0110;
	mem[761] = 4'b0101;
	mem[762] = 4'b0001;
	mem[763] = 4'b0000;
	mem[764] = 4'b0000;
	mem[765] = 4'b0000;
	mem[766] = 4'b0000;
	mem[767] = 4'b0000;
	mem[768] = 4'b0000;
	mem[769] = 4'b0000;
	mem[770] = 4'b0000;
	mem[771] = 4'b0000;
	mem[772] = 4'b0000;
	mem[773] = 4'b0000;
	mem[774] = 4'b0000;
	mem[775] = 4'b0000;
	mem[776] = 4'b0000;
	mem[777] = 4'b0001;
	mem[778] = 4'b0001;
	mem[779] = 4'b0001;
	mem[780] = 4'b0001;
	mem[781] = 4'b0001;
	mem[782] = 4'b0010;
	mem[783] = 4'b0011;
	mem[784] = 4'b0011;
	mem[785] = 4'b0011;
	mem[786] = 4'b0011;
	mem[787] = 4'b0011;
	mem[788] = 4'b0100;
	mem[789] = 4'b0100;
	mem[790] = 4'b0100;
	mem[791] = 4'b0101;
	mem[792] = 4'b0101;
	mem[793] = 4'b0101;
	mem[794] = 4'b0110;
	mem[795] = 4'b0110;
	mem[796] = 4'b0101;
	mem[797] = 4'b0101;
	mem[798] = 4'b0101;
	mem[799] = 4'b0110;
	mem[800] = 4'b0111;
	mem[801] = 4'b0111;
	mem[802] = 4'b0111;
	mem[803] = 4'b0111;
	mem[804] = 4'b0111;
	mem[805] = 4'b1000;
	mem[806] = 4'b1001;
	mem[807] = 4'b1010;
	mem[808] = 4'b1001;
	mem[809] = 4'b1001;
	mem[810] = 4'b1010;
	mem[811] = 4'b1011;
	mem[812] = 4'b1011;
	mem[813] = 4'b1011;
	mem[814] = 4'b1011;
	mem[815] = 4'b1011;
	mem[816] = 4'b1100;
	mem[817] = 4'b1100;
	mem[818] = 4'b1100;
	mem[819] = 4'b1100;
	mem[820] = 4'b1100;
	mem[821] = 4'b1101;
	mem[822] = 4'b1110;
	mem[823] = 4'b1110;
	mem[824] = 4'b1110;
	mem[825] = 4'b1110;
	mem[826] = 4'b1110;
	mem[827] = 4'b1111;
	mem[828] = 4'b1111;
	mem[829] = 4'b1111;
	mem[830] = 4'b1111;
	mem[831] = 4'b1111;
	mem[832] = 4'b1111;
	mem[833] = 4'b1111;
	mem[834] = 4'b1111;
	mem[835] = 4'b1111;
	mem[836] = 4'b1111;
	mem[837] = 4'b1110;
	mem[838] = 4'b0110;
	mem[839] = 4'b0001;
	mem[840] = 4'b0001;
	mem[841] = 4'b0001;
	mem[842] = 4'b0001;
	mem[843] = 4'b0010;
	mem[844] = 4'b0001;
	mem[845] = 4'b0001;
	mem[846] = 4'b0010;
	mem[847] = 4'b0010;
	mem[848] = 4'b0001;
	mem[849] = 4'b0010;
	mem[850] = 4'b0010;
	mem[851] = 4'b0010;
	mem[852] = 4'b0010;
	mem[853] = 4'b0010;
	mem[854] = 4'b0010;
	mem[855] = 4'b0010;
	mem[856] = 4'b0010;
	mem[857] = 4'b0010;
	mem[858] = 4'b0011;
	mem[859] = 4'b0011;
	mem[860] = 4'b0011;
	mem[861] = 4'b0011;
	mem[862] = 4'b0011;
	mem[863] = 4'b0011;
	mem[864] = 4'b0011;
	mem[865] = 4'b0011;
	mem[866] = 4'b0011;
	mem[867] = 4'b0100;
	mem[868] = 4'b0100;
	mem[869] = 4'b0100;
	mem[870] = 4'b0100;
	mem[871] = 4'b0100;
	mem[872] = 4'b0100;
	mem[873] = 4'b0100;
	mem[874] = 4'b0100;
	mem[875] = 4'b0100;
	mem[876] = 4'b0101;
	mem[877] = 4'b0101;
	mem[878] = 4'b0101;
	mem[879] = 4'b0101;
	mem[880] = 4'b0101;
	mem[881] = 4'b0101;
	mem[882] = 4'b0101;
	mem[883] = 4'b0101;
	mem[884] = 4'b0101;
	mem[885] = 4'b0101;
	mem[886] = 4'b0110;
	mem[887] = 4'b0110;
	mem[888] = 4'b0110;
	mem[889] = 4'b0110;
	mem[890] = 4'b0001;
	mem[891] = 4'b0000;
	mem[892] = 4'b0000;
	mem[893] = 4'b0000;
	mem[894] = 4'b0000;
	mem[895] = 4'b0000;
	mem[896] = 4'b0000;
	mem[897] = 4'b0000;
	mem[898] = 4'b0000;
	mem[899] = 4'b0000;
	mem[900] = 4'b0000;
	mem[901] = 4'b0000;
	mem[902] = 4'b0000;
	mem[903] = 4'b0000;
	mem[904] = 4'b0000;
	mem[905] = 4'b0001;
	mem[906] = 4'b0001;
	mem[907] = 4'b0001;
	mem[908] = 4'b0001;
	mem[909] = 4'b0001;
	mem[910] = 4'b0010;
	mem[911] = 4'b0011;
	mem[912] = 4'b0011;
	mem[913] = 4'b0011;
	mem[914] = 4'b0011;
	mem[915] = 4'b0011;
	mem[916] = 4'b0100;
	mem[917] = 4'b0100;
	mem[918] = 4'b0101;
	mem[919] = 4'b0101;
	mem[920] = 4'b0100;
	mem[921] = 4'b0101;
	mem[922] = 4'b0110;
	mem[923] = 4'b0110;
	mem[924] = 4'b0110;
	mem[925] = 4'b0110;
	mem[926] = 4'b0101;
	mem[927] = 4'b0110;
	mem[928] = 4'b0111;
	mem[929] = 4'b0111;
	mem[930] = 4'b0111;
	mem[931] = 4'b0111;
	mem[932] = 4'b0111;
	mem[933] = 4'b1001;
	mem[934] = 4'b1010;
	mem[935] = 4'b1001;
	mem[936] = 4'b1001;
	mem[937] = 4'b1001;
	mem[938] = 4'b1010;
	mem[939] = 4'b1011;
	mem[940] = 4'b1011;
	mem[941] = 4'b1011;
	mem[942] = 4'b1011;
	mem[943] = 4'b1011;
	mem[944] = 4'b1100;
	mem[945] = 4'b1100;
	mem[946] = 4'b1100;
	mem[947] = 4'b1100;
	mem[948] = 4'b1100;
	mem[949] = 4'b1101;
	mem[950] = 4'b1110;
	mem[951] = 4'b1110;
	mem[952] = 4'b1110;
	mem[953] = 4'b1110;
	mem[954] = 4'b1110;
	mem[955] = 4'b1111;
	mem[956] = 4'b1111;
	mem[957] = 4'b1111;
	mem[958] = 4'b1111;
	mem[959] = 4'b1111;
	mem[960] = 4'b1111;
	mem[961] = 4'b1111;
	mem[962] = 4'b1111;
	mem[963] = 4'b1111;
	mem[964] = 4'b1110;
	mem[965] = 4'b1101;
	mem[966] = 4'b0110;
	mem[967] = 4'b0001;
	mem[968] = 4'b0001;
	mem[969] = 4'b0001;
	mem[970] = 4'b0010;
	mem[971] = 4'b0001;
	mem[972] = 4'b0010;
	mem[973] = 4'b0010;
	mem[974] = 4'b0010;
	mem[975] = 4'b0010;
	mem[976] = 4'b0010;
	mem[977] = 4'b0010;
	mem[978] = 4'b0010;
	mem[979] = 4'b0010;
	mem[980] = 4'b0010;
	mem[981] = 4'b0010;
	mem[982] = 4'b0010;
	mem[983] = 4'b0010;
	mem[984] = 4'b0011;
	mem[985] = 4'b0011;
	mem[986] = 4'b0011;
	mem[987] = 4'b0011;
	mem[988] = 4'b0011;
	mem[989] = 4'b0011;
	mem[990] = 4'b0011;
	mem[991] = 4'b0011;
	mem[992] = 4'b0011;
	mem[993] = 4'b0100;
	mem[994] = 4'b0100;
	mem[995] = 4'b0100;
	mem[996] = 4'b0100;
	mem[997] = 4'b0100;
	mem[998] = 4'b0100;
	mem[999] = 4'b0100;
	mem[1000] = 4'b0100;
	mem[1001] = 4'b0100;
	mem[1002] = 4'b0101;
	mem[1003] = 4'b0101;
	mem[1004] = 4'b0101;
	mem[1005] = 4'b0101;
	mem[1006] = 4'b0101;
	mem[1007] = 4'b0101;
	mem[1008] = 4'b0101;
	mem[1009] = 4'b0101;
	mem[1010] = 4'b0101;
	mem[1011] = 4'b0110;
	mem[1012] = 4'b0110;
	mem[1013] = 4'b0110;
	mem[1014] = 4'b0110;
	mem[1015] = 4'b0110;
	mem[1016] = 4'b0110;
	mem[1017] = 4'b0110;
	mem[1018] = 4'b0001;
	mem[1019] = 4'b0000;
	mem[1020] = 4'b0000;
	mem[1021] = 4'b0000;
	mem[1022] = 4'b0000;
	mem[1023] = 4'b0000;
	mem[1024] = 4'b0000;
	mem[1025] = 4'b0000;
	mem[1026] = 4'b0000;
	mem[1027] = 4'b0000;
	mem[1028] = 4'b0000;
	mem[1029] = 4'b0000;
	mem[1030] = 4'b0000;
	mem[1031] = 4'b0000;
	mem[1032] = 4'b0000;
	mem[1033] = 4'b0001;
	mem[1034] = 4'b0001;
	mem[1035] = 4'b0001;
	mem[1036] = 4'b0001;
	mem[1037] = 4'b0001;
	mem[1038] = 4'b0010;
	mem[1039] = 4'b0011;
	mem[1040] = 4'b0011;
	mem[1041] = 4'b0011;
	mem[1042] = 4'b0011;
	mem[1043] = 4'b0100;
	mem[1044] = 4'b0101;
	mem[1045] = 4'b0101;
	mem[1046] = 4'b0101;
	mem[1047] = 4'b0100;
	mem[1048] = 4'b0100;
	mem[1049] = 4'b0101;
	mem[1050] = 4'b0110;
	mem[1051] = 4'b0110;
	mem[1052] = 4'b0110;
	mem[1053] = 4'b0110;
	mem[1054] = 4'b0110;
	mem[1055] = 4'b0111;
	mem[1056] = 4'b0111;
	mem[1057] = 4'b0111;
	mem[1058] = 4'b0111;
	mem[1059] = 4'b1000;
	mem[1060] = 4'b1000;
	mem[1061] = 4'b1001;
	mem[1062] = 4'b1001;
	mem[1063] = 4'b1001;
	mem[1064] = 4'b1001;
	mem[1065] = 4'b1001;
	mem[1066] = 4'b1010;
	mem[1067] = 4'b1011;
	mem[1068] = 4'b1011;
	mem[1069] = 4'b1011;
	mem[1070] = 4'b1011;
	mem[1071] = 4'b1011;
	mem[1072] = 4'b1100;
	mem[1073] = 4'b1100;
	mem[1074] = 4'b1100;
	mem[1075] = 4'b1100;
	mem[1076] = 4'b1100;
	mem[1077] = 4'b1101;
	mem[1078] = 4'b1110;
	mem[1079] = 4'b1110;
	mem[1080] = 4'b1110;
	mem[1081] = 4'b1110;
	mem[1082] = 4'b1110;
	mem[1083] = 4'b1111;
	mem[1084] = 4'b1111;
	mem[1085] = 4'b1111;
	mem[1086] = 4'b1111;
	mem[1087] = 4'b1111;
	mem[1088] = 4'b1111;
	mem[1089] = 4'b1111;
	mem[1090] = 4'b1111;
	mem[1091] = 4'b1110;
	mem[1092] = 4'b1101;
	mem[1093] = 4'b1110;
	mem[1094] = 4'b0111;
	mem[1095] = 4'b0010;
	mem[1096] = 4'b0001;
	mem[1097] = 4'b0001;
	mem[1098] = 4'b0010;
	mem[1099] = 4'b0010;
	mem[1100] = 4'b0010;
	mem[1101] = 4'b0010;
	mem[1102] = 4'b0010;
	mem[1103] = 4'b0011;
	mem[1104] = 4'b0011;
	mem[1105] = 4'b0010;
	mem[1106] = 4'b0010;
	mem[1107] = 4'b0010;
	mem[1108] = 4'b0010;
	mem[1109] = 4'b0011;
	mem[1110] = 4'b0011;
	mem[1111] = 4'b0011;
	mem[1112] = 4'b0011;
	mem[1113] = 4'b0011;
	mem[1114] = 4'b0011;
	mem[1115] = 4'b0011;
	mem[1116] = 4'b0011;
	mem[1117] = 4'b0011;
	mem[1118] = 4'b0100;
	mem[1119] = 4'b0100;
	mem[1120] = 4'b0100;
	mem[1121] = 4'b0100;
	mem[1122] = 4'b0100;
	mem[1123] = 4'b0100;
	mem[1124] = 4'b0100;
	mem[1125] = 4'b0100;
	mem[1126] = 4'b0100;
	mem[1127] = 4'b0101;
	mem[1128] = 4'b0101;
	mem[1129] = 4'b0101;
	mem[1130] = 4'b0101;
	mem[1131] = 4'b0101;
	mem[1132] = 4'b0101;
	mem[1133] = 4'b0101;
	mem[1134] = 4'b0101;
	mem[1135] = 4'b0101;
	mem[1136] = 4'b0101;
	mem[1137] = 4'b0110;
	mem[1138] = 4'b0110;
	mem[1139] = 4'b0110;
	mem[1140] = 4'b0110;
	mem[1141] = 4'b0110;
	mem[1142] = 4'b0110;
	mem[1143] = 4'b0110;
	mem[1144] = 4'b0110;
	mem[1145] = 4'b0110;
	mem[1146] = 4'b0001;
	mem[1147] = 4'b0000;
	mem[1148] = 4'b0000;
	mem[1149] = 4'b0000;
	mem[1150] = 4'b0000;
	mem[1151] = 4'b0000;
	mem[1152] = 4'b0000;
	mem[1153] = 4'b0000;
	mem[1154] = 4'b0000;
	mem[1155] = 4'b0000;
	mem[1156] = 4'b0000;
	mem[1157] = 4'b0000;
	mem[1158] = 4'b0000;
	mem[1159] = 4'b0000;
	mem[1160] = 4'b0000;
	mem[1161] = 4'b0001;
	mem[1162] = 4'b0001;
	mem[1163] = 4'b0001;
	mem[1164] = 4'b0001;
	mem[1165] = 4'b0001;
	mem[1166] = 4'b0010;
	mem[1167] = 4'b0011;
	mem[1168] = 4'b0011;
	mem[1169] = 4'b0011;
	mem[1170] = 4'b0100;
	mem[1171] = 4'b0011;
	mem[1172] = 4'b0100;
	mem[1173] = 4'b0101;
	mem[1174] = 4'b0101;
	mem[1175] = 4'b0100;
	mem[1176] = 4'b0100;
	mem[1177] = 4'b0101;
	mem[1178] = 4'b0110;
	mem[1179] = 4'b0110;
	mem[1180] = 4'b0110;
	mem[1181] = 4'b0110;
	mem[1182] = 4'b0110;
	mem[1183] = 4'b0111;
	mem[1184] = 4'b1000;
	mem[1185] = 4'b1000;
	mem[1186] = 4'b1000;
	mem[1187] = 4'b1000;
	mem[1188] = 4'b1000;
	mem[1189] = 4'b1001;
	mem[1190] = 4'b1001;
	mem[1191] = 4'b1001;
	mem[1192] = 4'b1001;
	mem[1193] = 4'b1001;
	mem[1194] = 4'b1010;
	mem[1195] = 4'b1011;
	mem[1196] = 4'b1011;
	mem[1197] = 4'b1011;
	mem[1198] = 4'b1011;
	mem[1199] = 4'b1011;
	mem[1200] = 4'b1100;
	mem[1201] = 4'b1100;
	mem[1202] = 4'b1100;
	mem[1203] = 4'b1100;
	mem[1204] = 4'b1100;
	mem[1205] = 4'b1101;
	mem[1206] = 4'b1110;
	mem[1207] = 4'b1110;
	mem[1208] = 4'b1110;
	mem[1209] = 4'b1110;
	mem[1210] = 4'b1110;
	mem[1211] = 4'b1111;
	mem[1212] = 4'b1111;
	mem[1213] = 4'b1111;
	mem[1214] = 4'b1111;
	mem[1215] = 4'b1111;
	mem[1216] = 4'b1111;
	mem[1217] = 4'b1111;
	mem[1218] = 4'b1111;
	mem[1219] = 4'b1101;
	mem[1220] = 4'b1110;
	mem[1221] = 4'b1111;
	mem[1222] = 4'b0111;
	mem[1223] = 4'b0001;
	mem[1224] = 4'b0010;
	mem[1225] = 4'b0010;
	mem[1226] = 4'b0010;
	mem[1227] = 4'b0011;
	mem[1228] = 4'b0010;
	mem[1229] = 4'b0010;
	mem[1230] = 4'b0011;
	mem[1231] = 4'b0011;
	mem[1232] = 4'b0011;
	mem[1233] = 4'b0010;
	mem[1234] = 4'b0010;
	mem[1235] = 4'b0011;
	mem[1236] = 4'b0011;
	mem[1237] = 4'b0011;
	mem[1238] = 4'b0011;
	mem[1239] = 4'b0011;
	mem[1240] = 4'b0011;
	mem[1241] = 4'b0011;
	mem[1242] = 4'b0011;
	mem[1243] = 4'b0011;
	mem[1244] = 4'b0100;
	mem[1245] = 4'b0100;
	mem[1246] = 4'b0100;
	mem[1247] = 4'b0100;
	mem[1248] = 4'b0100;
	mem[1249] = 4'b0100;
	mem[1250] = 4'b0100;
	mem[1251] = 4'b0100;
	mem[1252] = 4'b0100;
	mem[1253] = 4'b0101;
	mem[1254] = 4'b0101;
	mem[1255] = 4'b0101;
	mem[1256] = 4'b0101;
	mem[1257] = 4'b0101;
	mem[1258] = 4'b0101;
	mem[1259] = 4'b0101;
	mem[1260] = 4'b0101;
	mem[1261] = 4'b0101;
	mem[1262] = 4'b0110;
	mem[1263] = 4'b0110;
	mem[1264] = 4'b0110;
	mem[1265] = 4'b0110;
	mem[1266] = 4'b0110;
	mem[1267] = 4'b0110;
	mem[1268] = 4'b0110;
	mem[1269] = 4'b0110;
	mem[1270] = 4'b0110;
	mem[1271] = 4'b0111;
	mem[1272] = 4'b0111;
	mem[1273] = 4'b0110;
	mem[1274] = 4'b0001;
	mem[1275] = 4'b0000;
	mem[1276] = 4'b0000;
	mem[1277] = 4'b0000;
	mem[1278] = 4'b0000;
	mem[1279] = 4'b0000;
	mem[1280] = 4'b0000;
	mem[1281] = 4'b0000;
	mem[1282] = 4'b0000;
	mem[1283] = 4'b0000;
	mem[1284] = 4'b0000;
	mem[1285] = 4'b0000;
	mem[1286] = 4'b0000;
	mem[1287] = 4'b0000;
	mem[1288] = 4'b0000;
	mem[1289] = 4'b0001;
	mem[1290] = 4'b0001;
	mem[1291] = 4'b0001;
	mem[1292] = 4'b0001;
	mem[1293] = 4'b0001;
	mem[1294] = 4'b0010;
	mem[1295] = 4'b0011;
	mem[1296] = 4'b0011;
	mem[1297] = 4'b0100;
	mem[1298] = 4'b0011;
	mem[1299] = 4'b0011;
	mem[1300] = 4'b0100;
	mem[1301] = 4'b0100;
	mem[1302] = 4'b0100;
	mem[1303] = 4'b0100;
	mem[1304] = 4'b0100;
	mem[1305] = 4'b0101;
	mem[1306] = 4'b0110;
	mem[1307] = 4'b0101;
	mem[1308] = 4'b0110;
	mem[1309] = 4'b0110;
	mem[1310] = 4'b0110;
	mem[1311] = 4'b0111;
	mem[1312] = 4'b1000;
	mem[1313] = 4'b1000;
	mem[1314] = 4'b1000;
	mem[1315] = 4'b1000;
	mem[1316] = 4'b1000;
	mem[1317] = 4'b1001;
	mem[1318] = 4'b1001;
	mem[1319] = 4'b1001;
	mem[1320] = 4'b1001;
	mem[1321] = 4'b1001;
	mem[1322] = 4'b1010;
	mem[1323] = 4'b1011;
	mem[1324] = 4'b1011;
	mem[1325] = 4'b1011;
	mem[1326] = 4'b1011;
	mem[1327] = 4'b1011;
	mem[1328] = 4'b1100;
	mem[1329] = 4'b1100;
	mem[1330] = 4'b1100;
	mem[1331] = 4'b1100;
	mem[1332] = 4'b1100;
	mem[1333] = 4'b1101;
	mem[1334] = 4'b1110;
	mem[1335] = 4'b1110;
	mem[1336] = 4'b1110;
	mem[1337] = 4'b1110;
	mem[1338] = 4'b1110;
	mem[1339] = 4'b1111;
	mem[1340] = 4'b1111;
	mem[1341] = 4'b1111;
	mem[1342] = 4'b1111;
	mem[1343] = 4'b1111;
	mem[1344] = 4'b1111;
	mem[1345] = 4'b1111;
	mem[1346] = 4'b1110;
	mem[1347] = 4'b1101;
	mem[1348] = 4'b1110;
	mem[1349] = 4'b1111;
	mem[1350] = 4'b0111;
	mem[1351] = 4'b0010;
	mem[1352] = 4'b0010;
	mem[1353] = 4'b0010;
	mem[1354] = 4'b0010;
	mem[1355] = 4'b0011;
	mem[1356] = 4'b0011;
	mem[1357] = 4'b0010;
	mem[1358] = 4'b0010;
	mem[1359] = 4'b0011;
	mem[1360] = 4'b0011;
	mem[1361] = 4'b0011;
	mem[1362] = 4'b0011;
	mem[1363] = 4'b0011;
	mem[1364] = 4'b0011;
	mem[1365] = 4'b0011;
	mem[1366] = 4'b0011;
	mem[1367] = 4'b0011;
	mem[1368] = 4'b0011;
	mem[1369] = 4'b0100;
	mem[1370] = 4'b0100;
	mem[1371] = 4'b0100;
	mem[1372] = 4'b0100;
	mem[1373] = 4'b0100;
	mem[1374] = 4'b0100;
	mem[1375] = 4'b0100;
	mem[1376] = 4'b0100;
	mem[1377] = 4'b0100;
	mem[1378] = 4'b0101;
	mem[1379] = 4'b0101;
	mem[1380] = 4'b0101;
	mem[1381] = 4'b0101;
	mem[1382] = 4'b0101;
	mem[1383] = 4'b0101;
	mem[1384] = 4'b0101;
	mem[1385] = 4'b0101;
	mem[1386] = 4'b0101;
	mem[1387] = 4'b0110;
	mem[1388] = 4'b0110;
	mem[1389] = 4'b0110;
	mem[1390] = 4'b0110;
	mem[1391] = 4'b0110;
	mem[1392] = 4'b0110;
	mem[1393] = 4'b0110;
	mem[1394] = 4'b0110;
	mem[1395] = 4'b0110;
	mem[1396] = 4'b0110;
	mem[1397] = 4'b0111;
	mem[1398] = 4'b0111;
	mem[1399] = 4'b0111;
	mem[1400] = 4'b0111;
	mem[1401] = 4'b0111;
	mem[1402] = 4'b0001;
	mem[1403] = 4'b0000;
	mem[1404] = 4'b0000;
	mem[1405] = 4'b0000;
	mem[1406] = 4'b0000;
	mem[1407] = 4'b0000;
	mem[1408] = 4'b0000;
	mem[1409] = 4'b0000;
	mem[1410] = 4'b0000;
	mem[1411] = 4'b0000;
	mem[1412] = 4'b0000;
	mem[1413] = 4'b0000;
	mem[1414] = 4'b0000;
	mem[1415] = 4'b0000;
	mem[1416] = 4'b0000;
	mem[1417] = 4'b0001;
	mem[1418] = 4'b0001;
	mem[1419] = 4'b0001;
	mem[1420] = 4'b0001;
	mem[1421] = 4'b0001;
	mem[1422] = 4'b0010;
	mem[1423] = 4'b0011;
	mem[1424] = 4'b0011;
	mem[1425] = 4'b0100;
	mem[1426] = 4'b0011;
	mem[1427] = 4'b0011;
	mem[1428] = 4'b0100;
	mem[1429] = 4'b0100;
	mem[1430] = 4'b0100;
	mem[1431] = 4'b0100;
	mem[1432] = 4'b0100;
	mem[1433] = 4'b0101;
	mem[1434] = 4'b0101;
	mem[1435] = 4'b0101;
	mem[1436] = 4'b0110;
	mem[1437] = 4'b0110;
	mem[1438] = 4'b0110;
	mem[1439] = 4'b0111;
	mem[1440] = 4'b1000;
	mem[1441] = 4'b1000;
	mem[1442] = 4'b1000;
	mem[1443] = 4'b1000;
	mem[1444] = 4'b1000;
	mem[1445] = 4'b1001;
	mem[1446] = 4'b1001;
	mem[1447] = 4'b1001;
	mem[1448] = 4'b1001;
	mem[1449] = 4'b1001;
	mem[1450] = 4'b1010;
	mem[1451] = 4'b1011;
	mem[1452] = 4'b1011;
	mem[1453] = 4'b1011;
	mem[1454] = 4'b1011;
	mem[1455] = 4'b1011;
	mem[1456] = 4'b1100;
	mem[1457] = 4'b1100;
	mem[1458] = 4'b1100;
	mem[1459] = 4'b1100;
	mem[1460] = 4'b1100;
	mem[1461] = 4'b1101;
	mem[1462] = 4'b1110;
	mem[1463] = 4'b1110;
	mem[1464] = 4'b1110;
	mem[1465] = 4'b1110;
	mem[1466] = 4'b1110;
	mem[1467] = 4'b1111;
	mem[1468] = 4'b1111;
	mem[1469] = 4'b1111;
	mem[1470] = 4'b1111;
	mem[1471] = 4'b1111;
	mem[1472] = 4'b1111;
	mem[1473] = 4'b1111;
	mem[1474] = 4'b1110;
	mem[1475] = 4'b1101;
	mem[1476] = 4'b1110;
	mem[1477] = 4'b1111;
	mem[1478] = 4'b0111;
	mem[1479] = 4'b0010;
	mem[1480] = 4'b0010;
	mem[1481] = 4'b0010;
	mem[1482] = 4'b0010;
	mem[1483] = 4'b0011;
	mem[1484] = 4'b0011;
	mem[1485] = 4'b0011;
	mem[1486] = 4'b0011;
	mem[1487] = 4'b0011;
	mem[1488] = 4'b0011;
	mem[1489] = 4'b0011;
	mem[1490] = 4'b0011;
	mem[1491] = 4'b0011;
	mem[1492] = 4'b0011;
	mem[1493] = 4'b0011;
	mem[1494] = 4'b0011;
	mem[1495] = 4'b0100;
	mem[1496] = 4'b0100;
	mem[1497] = 4'b0100;
	mem[1498] = 4'b0100;
	mem[1499] = 4'b0100;
	mem[1500] = 4'b0100;
	mem[1501] = 4'b0100;
	mem[1502] = 4'b0100;
	mem[1503] = 4'b0100;
	mem[1504] = 4'b0101;
	mem[1505] = 4'b0101;
	mem[1506] = 4'b0101;
	mem[1507] = 4'b0101;
	mem[1508] = 4'b0101;
	mem[1509] = 4'b0101;
	mem[1510] = 4'b0101;
	mem[1511] = 4'b0101;
	mem[1512] = 4'b0101;
	mem[1513] = 4'b0110;
	mem[1514] = 4'b0110;
	mem[1515] = 4'b0110;
	mem[1516] = 4'b0110;
	mem[1517] = 4'b0110;
	mem[1518] = 4'b0110;
	mem[1519] = 4'b0110;
	mem[1520] = 4'b0110;
	mem[1521] = 4'b0110;
	mem[1522] = 4'b0111;
	mem[1523] = 4'b0111;
	mem[1524] = 4'b0111;
	mem[1525] = 4'b0111;
	mem[1526] = 4'b0111;
	mem[1527] = 4'b0111;
	mem[1528] = 4'b0111;
	mem[1529] = 4'b0111;
	mem[1530] = 4'b0001;
	mem[1531] = 4'b0000;
	mem[1532] = 4'b0000;
	mem[1533] = 4'b0000;
	mem[1534] = 4'b0000;
	mem[1535] = 4'b0000;
	mem[1536] = 4'b0000;
	mem[1537] = 4'b0000;
	mem[1538] = 4'b0000;
	mem[1539] = 4'b0000;
	mem[1540] = 4'b0000;
	mem[1541] = 4'b0000;
	mem[1542] = 4'b0000;
	mem[1543] = 4'b0000;
	mem[1544] = 4'b0000;
	mem[1545] = 4'b0001;
	mem[1546] = 4'b0001;
	mem[1547] = 4'b0001;
	mem[1548] = 4'b0001;
	mem[1549] = 4'b0001;
	mem[1550] = 4'b0010;
	mem[1551] = 4'b0010;
	mem[1552] = 4'b0010;
	mem[1553] = 4'b0011;
	mem[1554] = 4'b0010;
	mem[1555] = 4'b0010;
	mem[1556] = 4'b0100;
	mem[1557] = 4'b0100;
	mem[1558] = 4'b0100;
	mem[1559] = 4'b0100;
	mem[1560] = 4'b0100;
	mem[1561] = 4'b0100;
	mem[1562] = 4'b0101;
	mem[1563] = 4'b0101;
	mem[1564] = 4'b0101;
	mem[1565] = 4'b0110;
	mem[1566] = 4'b0101;
	mem[1567] = 4'b0110;
	mem[1568] = 4'b0111;
	mem[1569] = 4'b0111;
	mem[1570] = 4'b0111;
	mem[1571] = 4'b0111;
	mem[1572] = 4'b0111;
	mem[1573] = 4'b1000;
	mem[1574] = 4'b1000;
	mem[1575] = 4'b1000;
	mem[1576] = 4'b1000;
	mem[1577] = 4'b1000;
	mem[1578] = 4'b1001;
	mem[1579] = 4'b1010;
	mem[1580] = 4'b1010;
	mem[1581] = 4'b1010;
	mem[1582] = 4'b1010;
	mem[1583] = 4'b1010;
	mem[1584] = 4'b1011;
	mem[1585] = 4'b1011;
	mem[1586] = 4'b1011;
	mem[1587] = 4'b1011;
	mem[1588] = 4'b1011;
	mem[1589] = 4'b1100;
	mem[1590] = 4'b1101;
	mem[1591] = 4'b1101;
	mem[1592] = 4'b1101;
	mem[1593] = 4'b1101;
	mem[1594] = 4'b1101;
	mem[1595] = 4'b1101;
	mem[1596] = 4'b1101;
	mem[1597] = 4'b1101;
	mem[1598] = 4'b1101;
	mem[1599] = 4'b1101;
	mem[1600] = 4'b1101;
	mem[1601] = 4'b1110;
	mem[1602] = 4'b1110;
	mem[1603] = 4'b1100;
	mem[1604] = 4'b1100;
	mem[1605] = 4'b1101;
	mem[1606] = 4'b0111;
	mem[1607] = 4'b0010;
	mem[1608] = 4'b0010;
	mem[1609] = 4'b0010;
	mem[1610] = 4'b0010;
	mem[1611] = 4'b0011;
	mem[1612] = 4'b0011;
	mem[1613] = 4'b0010;
	mem[1614] = 4'b0011;
	mem[1615] = 4'b0011;
	mem[1616] = 4'b0011;
	mem[1617] = 4'b0011;
	mem[1618] = 4'b0011;
	mem[1619] = 4'b0011;
	mem[1620] = 4'b0011;
	mem[1621] = 4'b0011;
	mem[1622] = 4'b0011;
	mem[1623] = 4'b0011;
	mem[1624] = 4'b0100;
	mem[1625] = 4'b0100;
	mem[1626] = 4'b0100;
	mem[1627] = 4'b0100;
	mem[1628] = 4'b0100;
	mem[1629] = 4'b0100;
	mem[1630] = 4'b0100;
	mem[1631] = 4'b0100;
	mem[1632] = 4'b0100;
	mem[1633] = 4'b0100;
	mem[1634] = 4'b0101;
	mem[1635] = 4'b0101;
	mem[1636] = 4'b0101;
	mem[1637] = 4'b0101;
	mem[1638] = 4'b0101;
	mem[1639] = 4'b0101;
	mem[1640] = 4'b0101;
	mem[1641] = 4'b0101;
	mem[1642] = 4'b0101;
	mem[1643] = 4'b0101;
	mem[1644] = 4'b0110;
	mem[1645] = 4'b0110;
	mem[1646] = 4'b0110;
	mem[1647] = 4'b0110;
	mem[1648] = 4'b0110;
	mem[1649] = 4'b0110;
	mem[1650] = 4'b0110;
	mem[1651] = 4'b0110;
	mem[1652] = 4'b0110;
	mem[1653] = 4'b0110;
	mem[1654] = 4'b0111;
	mem[1655] = 4'b0111;
	mem[1656] = 4'b0111;
	mem[1657] = 4'b0111;
	mem[1658] = 4'b0001;
	mem[1659] = 4'b0000;
	mem[1660] = 4'b0000;
	mem[1661] = 4'b0000;
	mem[1662] = 4'b0000;
	mem[1663] = 4'b0000;
	mem[1664] = 4'b0000;
	mem[1665] = 4'b0000;
	mem[1666] = 4'b0000;
	mem[1667] = 4'b0000;
	mem[1668] = 4'b0000;
	mem[1669] = 4'b0000;
	mem[1670] = 4'b0000;
	mem[1671] = 4'b0000;
	mem[1672] = 4'b0000;
	mem[1673] = 4'b0000;
	mem[1674] = 4'b0000;
	mem[1675] = 4'b0000;
	mem[1676] = 4'b0000;
	mem[1677] = 4'b0000;
	mem[1678] = 4'b0000;
	mem[1679] = 4'b0000;
	mem[1680] = 4'b0000;
	mem[1681] = 4'b0001;
	mem[1682] = 4'b0000;
	mem[1683] = 4'b0000;
	mem[1684] = 4'b0000;
	mem[1685] = 4'b0000;
	mem[1686] = 4'b0000;
	mem[1687] = 4'b0000;
	mem[1688] = 4'b0000;
	mem[1689] = 4'b0001;
	mem[1690] = 4'b0000;
	mem[1691] = 4'b0001;
	mem[1692] = 4'b0001;
	mem[1693] = 4'b0001;
	mem[1694] = 4'b0000;
	mem[1695] = 4'b0000;
	mem[1696] = 4'b0000;
	mem[1697] = 4'b0000;
	mem[1698] = 4'b0000;
	mem[1699] = 4'b0000;
	mem[1700] = 4'b0000;
	mem[1701] = 4'b0000;
	mem[1702] = 4'b0000;
	mem[1703] = 4'b0000;
	mem[1704] = 4'b0000;
	mem[1705] = 4'b0000;
	mem[1706] = 4'b0000;
	mem[1707] = 4'b0001;
	mem[1708] = 4'b0001;
	mem[1709] = 4'b0001;
	mem[1710] = 4'b0001;
	mem[1711] = 4'b0001;
	mem[1712] = 4'b0001;
	mem[1713] = 4'b0001;
	mem[1714] = 4'b0001;
	mem[1715] = 4'b0001;
	mem[1716] = 4'b0001;
	mem[1717] = 4'b0001;
	mem[1718] = 4'b0001;
	mem[1719] = 4'b0001;
	mem[1720] = 4'b0001;
	mem[1721] = 4'b0001;
	mem[1722] = 4'b0001;
	mem[1723] = 4'b0001;
	mem[1724] = 4'b0001;
	mem[1725] = 4'b0001;
	mem[1726] = 4'b0001;
	mem[1727] = 4'b0001;
	mem[1728] = 4'b0001;
	mem[1729] = 4'b0010;
	mem[1730] = 4'b0001;
	mem[1731] = 4'b0010;
	mem[1732] = 4'b0001;
	mem[1733] = 4'b0001;
	mem[1734] = 4'b0001;
	mem[1735] = 4'b0000;
	mem[1736] = 4'b0000;
	mem[1737] = 4'b0000;
	mem[1738] = 4'b0001;
	mem[1739] = 4'b0001;
	mem[1740] = 4'b0000;
	mem[1741] = 4'b0000;
	mem[1742] = 4'b0000;
	mem[1743] = 4'b0000;
	mem[1744] = 4'b0000;
	mem[1745] = 4'b0000;
	mem[1746] = 4'b0000;
	mem[1747] = 4'b0000;
	mem[1748] = 4'b0000;
	mem[1749] = 4'b0000;
	mem[1750] = 4'b0000;
	mem[1751] = 4'b0000;
	mem[1752] = 4'b0000;
	mem[1753] = 4'b0000;
	mem[1754] = 4'b0000;
	mem[1755] = 4'b0000;
	mem[1756] = 4'b0000;
	mem[1757] = 4'b0000;
	mem[1758] = 4'b0000;
	mem[1759] = 4'b0000;
	mem[1760] = 4'b0000;
	mem[1761] = 4'b0000;
	mem[1762] = 4'b0000;
	mem[1763] = 4'b0000;
	mem[1764] = 4'b0000;
	mem[1765] = 4'b0000;
	mem[1766] = 4'b0000;
	mem[1767] = 4'b0000;
	mem[1768] = 4'b0000;
	mem[1769] = 4'b0000;
	mem[1770] = 4'b0000;
	mem[1771] = 4'b0000;
	mem[1772] = 4'b0000;
	mem[1773] = 4'b0000;
	mem[1774] = 4'b0000;
	mem[1775] = 4'b0000;
	mem[1776] = 4'b0000;
	mem[1777] = 4'b0000;
	mem[1778] = 4'b0000;
	mem[1779] = 4'b0000;
	mem[1780] = 4'b0000;
	mem[1781] = 4'b0000;
	mem[1782] = 4'b0000;
	mem[1783] = 4'b0000;
	mem[1784] = 4'b0000;
	mem[1785] = 4'b0000;
	mem[1786] = 4'b0000;
	mem[1787] = 4'b0000;
	mem[1788] = 4'b0000;
	mem[1789] = 4'b0000;
	mem[1790] = 4'b0000;
	mem[1791] = 4'b0000;
	mem[1792] = 4'b0000;
	mem[1793] = 4'b0000;
	mem[1794] = 4'b0000;
	mem[1795] = 4'b0000;
	mem[1796] = 4'b0000;
	mem[1797] = 4'b0000;
	mem[1798] = 4'b0000;
	mem[1799] = 4'b0000;
	mem[1800] = 4'b0000;
	mem[1801] = 4'b0000;
	mem[1802] = 4'b0000;
	mem[1803] = 4'b0000;
	mem[1804] = 4'b0000;
	mem[1805] = 4'b0000;
	mem[1806] = 4'b0000;
	mem[1807] = 4'b0000;
	mem[1808] = 4'b0000;
	mem[1809] = 4'b0000;
	mem[1810] = 4'b0001;
	mem[1811] = 4'b0000;
	mem[1812] = 4'b0000;
	mem[1813] = 4'b0000;
	mem[1814] = 4'b0000;
	mem[1815] = 4'b0000;
	mem[1816] = 4'b0000;
	mem[1817] = 4'b0000;
	mem[1818] = 4'b0000;
	mem[1819] = 4'b0000;
	mem[1820] = 4'b0000;
	mem[1821] = 4'b0001;
	mem[1822] = 4'b0000;
	mem[1823] = 4'b0000;
	mem[1824] = 4'b0000;
	mem[1825] = 4'b0000;
	mem[1826] = 4'b0000;
	mem[1827] = 4'b0000;
	mem[1828] = 4'b0000;
	mem[1829] = 4'b0000;
	mem[1830] = 4'b0000;
	mem[1831] = 4'b0000;
	mem[1832] = 4'b0000;
	mem[1833] = 4'b0000;
	mem[1834] = 4'b0000;
	mem[1835] = 4'b0000;
	mem[1836] = 4'b0000;
	mem[1837] = 4'b0000;
	mem[1838] = 4'b0000;
	mem[1839] = 4'b0000;
	mem[1840] = 4'b0000;
	mem[1841] = 4'b0000;
	mem[1842] = 4'b0000;
	mem[1843] = 4'b0000;
	mem[1844] = 4'b0000;
	mem[1845] = 4'b0000;
	mem[1846] = 4'b0000;
	mem[1847] = 4'b0000;
	mem[1848] = 4'b0000;
	mem[1849] = 4'b0000;
	mem[1850] = 4'b0000;
	mem[1851] = 4'b0000;
	mem[1852] = 4'b0000;
	mem[1853] = 4'b0000;
	mem[1854] = 4'b0000;
	mem[1855] = 4'b0000;
	mem[1856] = 4'b0000;
	mem[1857] = 4'b0001;
	mem[1858] = 4'b0000;
	mem[1859] = 4'b0000;
	mem[1860] = 4'b0000;
	mem[1861] = 4'b0000;
	mem[1862] = 4'b0000;
	mem[1863] = 4'b0000;
	mem[1864] = 4'b0000;
	mem[1865] = 4'b0001;
	mem[1866] = 4'b0001;
	mem[1867] = 4'b0000;
	mem[1868] = 4'b0000;
	mem[1869] = 4'b0000;
	mem[1870] = 4'b0000;
	mem[1871] = 4'b0000;
	mem[1872] = 4'b0000;
	mem[1873] = 4'b0000;
	mem[1874] = 4'b0000;
	mem[1875] = 4'b0000;
	mem[1876] = 4'b0000;
	mem[1877] = 4'b0000;
	mem[1878] = 4'b0000;
	mem[1879] = 4'b0000;
	mem[1880] = 4'b0000;
	mem[1881] = 4'b0000;
	mem[1882] = 4'b0000;
	mem[1883] = 4'b0000;
	mem[1884] = 4'b0000;
	mem[1885] = 4'b0000;
	mem[1886] = 4'b0000;
	mem[1887] = 4'b0000;
	mem[1888] = 4'b0000;
	mem[1889] = 4'b0000;
	mem[1890] = 4'b0000;
	mem[1891] = 4'b0000;
	mem[1892] = 4'b0000;
	mem[1893] = 4'b0000;
	mem[1894] = 4'b0000;
	mem[1895] = 4'b0000;
	mem[1896] = 4'b0000;
	mem[1897] = 4'b0000;
	mem[1898] = 4'b0000;
	mem[1899] = 4'b0000;
	mem[1900] = 4'b0000;
	mem[1901] = 4'b0000;
	mem[1902] = 4'b0000;
	mem[1903] = 4'b0000;
	mem[1904] = 4'b0000;
	mem[1905] = 4'b0000;
	mem[1906] = 4'b0000;
	mem[1907] = 4'b0000;
	mem[1908] = 4'b0000;
	mem[1909] = 4'b0000;
	mem[1910] = 4'b0000;
	mem[1911] = 4'b0000;
	mem[1912] = 4'b0000;
	mem[1913] = 4'b0000;
	mem[1914] = 4'b0000;
	mem[1915] = 4'b0000;
	mem[1916] = 4'b0000;
	mem[1917] = 4'b0000;
	mem[1918] = 4'b0000;
	mem[1919] = 4'b0000;
	mem[1920] = 4'b0000;
	mem[1921] = 4'b0000;
	mem[1922] = 4'b0000;
	mem[1923] = 4'b0000;
	mem[1924] = 4'b0000;
	mem[1925] = 4'b0000;
	mem[1926] = 4'b0000;
	mem[1927] = 4'b0000;
	mem[1928] = 4'b0000;
	mem[1929] = 4'b0000;
	mem[1930] = 4'b0000;
	mem[1931] = 4'b0000;
	mem[1932] = 4'b0000;
	mem[1933] = 4'b0000;
	mem[1934] = 4'b0000;
	mem[1935] = 4'b0000;
	mem[1936] = 4'b0000;
	mem[1937] = 4'b0000;
	mem[1938] = 4'b0000;
	mem[1939] = 4'b0000;
	mem[1940] = 4'b0000;
	mem[1941] = 4'b0000;
	mem[1942] = 4'b0000;
	mem[1943] = 4'b0000;
	mem[1944] = 4'b0000;
	mem[1945] = 4'b0000;
	mem[1946] = 4'b0000;
	mem[1947] = 4'b0000;
	mem[1948] = 4'b0001;
	mem[1949] = 4'b0000;
	mem[1950] = 4'b0000;
	mem[1951] = 4'b0000;
	mem[1952] = 4'b0000;
	mem[1953] = 4'b0000;
	mem[1954] = 4'b0000;
	mem[1955] = 4'b0000;
	mem[1956] = 4'b0000;
	mem[1957] = 4'b0000;
	mem[1958] = 4'b0000;
	mem[1959] = 4'b0000;
	mem[1960] = 4'b0000;
	mem[1961] = 4'b0000;
	mem[1962] = 4'b0000;
	mem[1963] = 4'b0000;
	mem[1964] = 4'b0000;
	mem[1965] = 4'b0000;
	mem[1966] = 4'b0000;
	mem[1967] = 4'b0000;
	mem[1968] = 4'b0000;
	mem[1969] = 4'b0000;
	mem[1970] = 4'b0000;
	mem[1971] = 4'b0000;
	mem[1972] = 4'b0000;
	mem[1973] = 4'b0000;
	mem[1974] = 4'b0000;
	mem[1975] = 4'b0000;
	mem[1976] = 4'b0000;
	mem[1977] = 4'b0000;
	mem[1978] = 4'b0000;
	mem[1979] = 4'b0000;
	mem[1980] = 4'b0000;
	mem[1981] = 4'b0000;
	mem[1982] = 4'b0001;
	mem[1983] = 4'b0001;
	mem[1984] = 4'b0001;
	mem[1985] = 4'b0000;
	mem[1986] = 4'b0000;
	mem[1987] = 4'b0000;
	mem[1988] = 4'b0000;
	mem[1989] = 4'b0000;
	mem[1990] = 4'b0001;
	mem[1991] = 4'b0001;
	mem[1992] = 4'b0001;
	mem[1993] = 4'b0001;
	mem[1994] = 4'b0000;
	mem[1995] = 4'b0000;
	mem[1996] = 4'b0000;
	mem[1997] = 4'b0000;
	mem[1998] = 4'b0000;
	mem[1999] = 4'b0000;
	mem[2000] = 4'b0000;
	mem[2001] = 4'b0000;
	mem[2002] = 4'b0000;
	mem[2003] = 4'b0000;
	mem[2004] = 4'b0000;
	mem[2005] = 4'b0000;
	mem[2006] = 4'b0000;
	mem[2007] = 4'b0000;
	mem[2008] = 4'b0000;
	mem[2009] = 4'b0000;
	mem[2010] = 4'b0000;
	mem[2011] = 4'b0000;
	mem[2012] = 4'b0000;
	mem[2013] = 4'b0000;
	mem[2014] = 4'b0000;
	mem[2015] = 4'b0000;
	mem[2016] = 4'b0000;
	mem[2017] = 4'b0000;
	mem[2018] = 4'b0000;
	mem[2019] = 4'b0000;
	mem[2020] = 4'b0000;
	mem[2021] = 4'b0000;
	mem[2022] = 4'b0000;
	mem[2023] = 4'b0000;
	mem[2024] = 4'b0000;
	mem[2025] = 4'b0000;
	mem[2026] = 4'b0000;
	mem[2027] = 4'b0000;
	mem[2028] = 4'b0000;
	mem[2029] = 4'b0000;
	mem[2030] = 4'b0000;
	mem[2031] = 4'b0000;
	mem[2032] = 4'b0000;
	mem[2033] = 4'b0000;
	mem[2034] = 4'b0000;
	mem[2035] = 4'b0000;
	mem[2036] = 4'b0000;
	mem[2037] = 4'b0000;
	mem[2038] = 4'b0000;
	mem[2039] = 4'b0000;
	mem[2040] = 4'b0000;
	mem[2041] = 4'b0000;
	mem[2042] = 4'b0000;
	mem[2043] = 4'b0000;
	mem[2044] = 4'b0000;
	mem[2045] = 4'b0000;
	mem[2046] = 4'b0000;
	mem[2047] = 4'b0000;
	mem[2048] = 4'b0000;
	mem[2049] = 4'b0000;
	mem[2050] = 4'b0000;
	mem[2051] = 4'b0000;
	mem[2052] = 4'b0000;
	mem[2053] = 4'b0000;
	mem[2054] = 4'b0000;
	mem[2055] = 4'b0000;
	mem[2056] = 4'b0000;
	mem[2057] = 4'b0000;
	mem[2058] = 4'b0000;
	mem[2059] = 4'b0000;
	mem[2060] = 4'b0000;
	mem[2061] = 4'b0000;
	mem[2062] = 4'b0000;
	mem[2063] = 4'b0000;
	mem[2064] = 4'b0000;
	mem[2065] = 4'b0000;
	mem[2066] = 4'b0000;
	mem[2067] = 4'b0000;
	mem[2068] = 4'b0000;
	mem[2069] = 4'b0000;
	mem[2070] = 4'b0000;
	mem[2071] = 4'b0000;
	mem[2072] = 4'b0000;
	mem[2073] = 4'b0000;
	mem[2074] = 4'b0000;
	mem[2075] = 4'b0000;
	mem[2076] = 4'b0001;
	mem[2077] = 4'b0000;
	mem[2078] = 4'b0000;
	mem[2079] = 4'b0000;
	mem[2080] = 4'b0000;
	mem[2081] = 4'b0000;
	mem[2082] = 4'b0000;
	mem[2083] = 4'b0000;
	mem[2084] = 4'b0000;
	mem[2085] = 4'b0000;
	mem[2086] = 4'b0000;
	mem[2087] = 4'b0000;
	mem[2088] = 4'b0000;
	mem[2089] = 4'b0000;
	mem[2090] = 4'b0000;
	mem[2091] = 4'b0000;
	mem[2092] = 4'b0000;
	mem[2093] = 4'b0000;
	mem[2094] = 4'b0000;
	mem[2095] = 4'b0000;
	mem[2096] = 4'b0000;
	mem[2097] = 4'b0000;
	mem[2098] = 4'b0000;
	mem[2099] = 4'b0000;
	mem[2100] = 4'b0000;
	mem[2101] = 4'b0000;
	mem[2102] = 4'b0000;
	mem[2103] = 4'b0000;
	mem[2104] = 4'b0000;
	mem[2105] = 4'b0000;
	mem[2106] = 4'b0000;
	mem[2107] = 4'b0000;
	mem[2108] = 4'b0000;
	mem[2109] = 4'b0000;
	mem[2110] = 4'b0001;
	mem[2111] = 4'b0000;
	mem[2112] = 4'b0000;
	mem[2113] = 4'b0000;
	mem[2114] = 4'b0000;
	mem[2115] = 4'b0000;
	mem[2116] = 4'b0000;
	mem[2117] = 4'b0000;
	mem[2118] = 4'b0000;
	mem[2119] = 4'b0000;
	mem[2120] = 4'b0000;
	mem[2121] = 4'b0000;
	mem[2122] = 4'b0000;
	mem[2123] = 4'b0000;
	mem[2124] = 4'b0000;
	mem[2125] = 4'b0000;
	mem[2126] = 4'b0000;
	mem[2127] = 4'b0000;
	mem[2128] = 4'b0000;
	mem[2129] = 4'b0000;
	mem[2130] = 4'b0000;
	mem[2131] = 4'b0000;
	mem[2132] = 4'b0000;
	mem[2133] = 4'b0000;
	mem[2134] = 4'b0000;
	mem[2135] = 4'b0000;
	mem[2136] = 4'b0000;
	mem[2137] = 4'b0000;
	mem[2138] = 4'b0000;
	mem[2139] = 4'b0000;
	mem[2140] = 4'b0000;
	mem[2141] = 4'b0000;
	mem[2142] = 4'b0000;
	mem[2143] = 4'b0000;
	mem[2144] = 4'b0000;
	mem[2145] = 4'b0000;
	mem[2146] = 4'b0000;
	mem[2147] = 4'b0000;
	mem[2148] = 4'b0000;
	mem[2149] = 4'b0000;
	mem[2150] = 4'b0000;
	mem[2151] = 4'b0000;
	mem[2152] = 4'b0000;
	mem[2153] = 4'b0000;
	mem[2154] = 4'b0000;
	mem[2155] = 4'b0000;
	mem[2156] = 4'b0000;
	mem[2157] = 4'b0000;
	mem[2158] = 4'b0000;
	mem[2159] = 4'b0000;
	mem[2160] = 4'b0000;
	mem[2161] = 4'b0000;
	mem[2162] = 4'b0000;
	mem[2163] = 4'b0000;
	mem[2164] = 4'b0000;
	mem[2165] = 4'b0000;
	mem[2166] = 4'b0000;
	mem[2167] = 4'b0000;
	mem[2168] = 4'b0000;
	mem[2169] = 4'b0000;
	mem[2170] = 4'b0000;
	mem[2171] = 4'b0000;
	mem[2172] = 4'b0000;
	mem[2173] = 4'b0000;
	mem[2174] = 4'b0000;
	mem[2175] = 4'b0000;
	mem[2176] = 4'b0000;
	mem[2177] = 4'b0000;
	mem[2178] = 4'b0000;
	mem[2179] = 4'b0000;
	mem[2180] = 4'b0000;
	mem[2181] = 4'b0000;
	mem[2182] = 4'b0000;
	mem[2183] = 4'b0000;
	mem[2184] = 4'b0000;
	mem[2185] = 4'b0000;
	mem[2186] = 4'b0000;
	mem[2187] = 4'b0000;
	mem[2188] = 4'b0000;
	mem[2189] = 4'b0000;
	mem[2190] = 4'b0000;
	mem[2191] = 4'b0000;
	mem[2192] = 4'b0000;
	mem[2193] = 4'b0000;
	mem[2194] = 4'b0000;
	mem[2195] = 4'b0000;
	mem[2196] = 4'b0000;
	mem[2197] = 4'b0000;
	mem[2198] = 4'b0000;
	mem[2199] = 4'b0000;
	mem[2200] = 4'b0000;
	mem[2201] = 4'b0000;
	mem[2202] = 4'b0000;
	mem[2203] = 4'b0001;
	mem[2204] = 4'b0000;
	mem[2205] = 4'b0000;
	mem[2206] = 4'b0000;
	mem[2207] = 4'b0000;
	mem[2208] = 4'b0000;
	mem[2209] = 4'b0000;
	mem[2210] = 4'b0000;
	mem[2211] = 4'b0000;
	mem[2212] = 4'b0000;
	mem[2213] = 4'b0000;
	mem[2214] = 4'b0000;
	mem[2215] = 4'b0000;
	mem[2216] = 4'b0000;
	mem[2217] = 4'b0000;
	mem[2218] = 4'b0000;
	mem[2219] = 4'b0000;
	mem[2220] = 4'b0000;
	mem[2221] = 4'b0000;
	mem[2222] = 4'b0000;
	mem[2223] = 4'b0000;
	mem[2224] = 4'b0000;
	mem[2225] = 4'b0000;
	mem[2226] = 4'b0000;
	mem[2227] = 4'b0000;
	mem[2228] = 4'b0000;
	mem[2229] = 4'b0000;
	mem[2230] = 4'b0000;
	mem[2231] = 4'b0000;
	mem[2232] = 4'b0000;
	mem[2233] = 4'b0000;
	mem[2234] = 4'b0000;
	mem[2235] = 4'b0000;
	mem[2236] = 4'b0000;
	mem[2237] = 4'b0000;
	mem[2238] = 4'b0001;
	mem[2239] = 4'b0000;
	mem[2240] = 4'b0000;
	mem[2241] = 4'b0000;
	mem[2242] = 4'b0000;
	mem[2243] = 4'b0000;
	mem[2244] = 4'b0000;
	mem[2245] = 4'b0000;
	mem[2246] = 4'b0000;
	mem[2247] = 4'b0000;
	mem[2248] = 4'b0000;
	mem[2249] = 4'b0000;
	mem[2250] = 4'b0000;
	mem[2251] = 4'b0000;
	mem[2252] = 4'b0000;
	mem[2253] = 4'b0000;
	mem[2254] = 4'b0000;
	mem[2255] = 4'b0000;
	mem[2256] = 4'b0000;
	mem[2257] = 4'b0000;
	mem[2258] = 4'b0000;
	mem[2259] = 4'b0000;
	mem[2260] = 4'b0000;
	mem[2261] = 4'b0000;
	mem[2262] = 4'b0000;
	mem[2263] = 4'b0000;
	mem[2264] = 4'b0000;
	mem[2265] = 4'b0000;
	mem[2266] = 4'b0000;
	mem[2267] = 4'b0000;
	mem[2268] = 4'b0000;
	mem[2269] = 4'b0000;
	mem[2270] = 4'b0000;
	mem[2271] = 4'b0000;
	mem[2272] = 4'b0000;
	mem[2273] = 4'b0000;
	mem[2274] = 4'b0000;
	mem[2275] = 4'b0000;
	mem[2276] = 4'b0000;
	mem[2277] = 4'b0000;
	mem[2278] = 4'b0000;
	mem[2279] = 4'b0000;
	mem[2280] = 4'b0000;
	mem[2281] = 4'b0000;
	mem[2282] = 4'b0000;
	mem[2283] = 4'b0000;
	mem[2284] = 4'b0000;
	mem[2285] = 4'b0000;
	mem[2286] = 4'b0000;
	mem[2287] = 4'b0000;
	mem[2288] = 4'b0000;
	mem[2289] = 4'b0000;
	mem[2290] = 4'b0000;
	mem[2291] = 4'b0000;
	mem[2292] = 4'b0000;
	mem[2293] = 4'b0000;
	mem[2294] = 4'b0000;
	mem[2295] = 4'b0000;
	mem[2296] = 4'b0000;
	mem[2297] = 4'b0000;
	mem[2298] = 4'b0000;
	mem[2299] = 4'b0000;
	mem[2300] = 4'b0000;
	mem[2301] = 4'b0000;
	mem[2302] = 4'b0000;
	mem[2303] = 4'b0000;
	mem[2304] = 4'b0000;
	mem[2305] = 4'b0000;
	mem[2306] = 4'b0000;
	mem[2307] = 4'b0000;
	mem[2308] = 4'b0000;
	mem[2309] = 4'b0000;
	mem[2310] = 4'b0000;
	mem[2311] = 4'b0000;
	mem[2312] = 4'b0000;
	mem[2313] = 4'b0000;
	mem[2314] = 4'b0000;
	mem[2315] = 4'b0000;
	mem[2316] = 4'b0000;
	mem[2317] = 4'b0000;
	mem[2318] = 4'b0000;
	mem[2319] = 4'b0000;
	mem[2320] = 4'b0000;
	mem[2321] = 4'b0000;
	mem[2322] = 4'b0000;
	mem[2323] = 4'b0000;
	mem[2324] = 4'b0000;
	mem[2325] = 4'b0000;
	mem[2326] = 4'b0000;
	mem[2327] = 4'b0000;
	mem[2328] = 4'b0000;
	mem[2329] = 4'b0000;
	mem[2330] = 4'b0001;
	mem[2331] = 4'b0001;
	mem[2332] = 4'b0000;
	mem[2333] = 4'b0000;
	mem[2334] = 4'b0000;
	mem[2335] = 4'b0000;
	mem[2336] = 4'b0000;
	mem[2337] = 4'b0000;
	mem[2338] = 4'b0000;
	mem[2339] = 4'b0000;
	mem[2340] = 4'b0000;
	mem[2341] = 4'b0000;
	mem[2342] = 4'b0000;
	mem[2343] = 4'b0000;
	mem[2344] = 4'b0000;
	mem[2345] = 4'b0000;
	mem[2346] = 4'b0000;
	mem[2347] = 4'b0000;
	mem[2348] = 4'b0000;
	mem[2349] = 4'b0000;
	mem[2350] = 4'b0000;
	mem[2351] = 4'b0000;
	mem[2352] = 4'b0000;
	mem[2353] = 4'b0000;
	mem[2354] = 4'b0000;
	mem[2355] = 4'b0000;
	mem[2356] = 4'b0000;
	mem[2357] = 4'b0000;
	mem[2358] = 4'b0000;
	mem[2359] = 4'b0000;
	mem[2360] = 4'b0000;
	mem[2361] = 4'b0000;
	mem[2362] = 4'b0000;
	mem[2363] = 4'b0000;
	mem[2364] = 4'b0000;
	mem[2365] = 4'b0000;
	mem[2366] = 4'b0000;
	mem[2367] = 4'b0000;
	mem[2368] = 4'b0000;
	mem[2369] = 4'b0000;
	mem[2370] = 4'b0000;
	mem[2371] = 4'b0000;
	mem[2372] = 4'b0001;
	mem[2373] = 4'b0000;
	mem[2374] = 4'b0000;
	mem[2375] = 4'b0000;
	mem[2376] = 4'b0000;
	mem[2377] = 4'b0000;
	mem[2378] = 4'b0000;
	mem[2379] = 4'b0000;
	mem[2380] = 4'b0000;
	mem[2381] = 4'b0000;
	mem[2382] = 4'b0000;
	mem[2383] = 4'b0000;
	mem[2384] = 4'b0000;
	mem[2385] = 4'b0000;
	mem[2386] = 4'b0000;
	mem[2387] = 4'b0000;
	mem[2388] = 4'b0000;
	mem[2389] = 4'b0000;
	mem[2390] = 4'b0000;
	mem[2391] = 4'b0000;
	mem[2392] = 4'b0000;
	mem[2393] = 4'b0000;
	mem[2394] = 4'b0000;
	mem[2395] = 4'b0000;
	mem[2396] = 4'b0000;
	mem[2397] = 4'b0000;
	mem[2398] = 4'b0000;
	mem[2399] = 4'b0000;
	mem[2400] = 4'b0000;
	mem[2401] = 4'b0000;
	mem[2402] = 4'b0000;
	mem[2403] = 4'b0000;
	mem[2404] = 4'b0000;
	mem[2405] = 4'b0000;
	mem[2406] = 4'b0000;
	mem[2407] = 4'b0000;
	mem[2408] = 4'b0000;
	mem[2409] = 4'b0000;
	mem[2410] = 4'b0000;
	mem[2411] = 4'b0000;
	mem[2412] = 4'b0000;
	mem[2413] = 4'b0000;
	mem[2414] = 4'b0000;
	mem[2415] = 4'b0000;
	mem[2416] = 4'b0000;
	mem[2417] = 4'b0000;
	mem[2418] = 4'b0000;
	mem[2419] = 4'b0000;
	mem[2420] = 4'b0000;
	mem[2421] = 4'b0000;
	mem[2422] = 4'b0000;
	mem[2423] = 4'b0000;
	mem[2424] = 4'b0000;
	mem[2425] = 4'b0000;
	mem[2426] = 4'b0000;
	mem[2427] = 4'b0000;
	mem[2428] = 4'b0000;
	mem[2429] = 4'b0000;
	mem[2430] = 4'b0000;
	mem[2431] = 4'b0000;
	mem[2432] = 4'b0000;
	mem[2433] = 4'b0000;
	mem[2434] = 4'b0000;
	mem[2435] = 4'b0000;
	mem[2436] = 4'b0000;
	mem[2437] = 4'b0000;
	mem[2438] = 4'b0000;
	mem[2439] = 4'b0000;
	mem[2440] = 4'b0000;
	mem[2441] = 4'b0000;
	mem[2442] = 4'b0000;
	mem[2443] = 4'b0000;
	mem[2444] = 4'b0000;
	mem[2445] = 4'b0000;
	mem[2446] = 4'b0000;
	mem[2447] = 4'b0000;
	mem[2448] = 4'b0000;
	mem[2449] = 4'b0000;
	mem[2450] = 4'b0000;
	mem[2451] = 4'b0000;
	mem[2452] = 4'b0000;
	mem[2453] = 4'b0000;
	mem[2454] = 4'b0000;
	mem[2455] = 4'b0000;
	mem[2456] = 4'b0000;
	mem[2457] = 4'b0001;
	mem[2458] = 4'b0001;
	mem[2459] = 4'b0000;
	mem[2460] = 4'b0000;
	mem[2461] = 4'b0000;
	mem[2462] = 4'b0000;
	mem[2463] = 4'b0000;
	mem[2464] = 4'b0000;
	mem[2465] = 4'b0000;
	mem[2466] = 4'b0000;
	mem[2467] = 4'b0000;
	mem[2468] = 4'b0000;
	mem[2469] = 4'b0000;
	mem[2470] = 4'b0000;
	mem[2471] = 4'b0000;
	mem[2472] = 4'b0000;
	mem[2473] = 4'b0000;
	mem[2474] = 4'b0000;
	mem[2475] = 4'b0000;
	mem[2476] = 4'b0000;
	mem[2477] = 4'b0000;
	mem[2478] = 4'b0000;
	mem[2479] = 4'b0000;
	mem[2480] = 4'b0000;
	mem[2481] = 4'b0000;
	mem[2482] = 4'b0000;
	mem[2483] = 4'b0000;
	mem[2484] = 4'b0000;
	mem[2485] = 4'b0000;
	mem[2486] = 4'b0000;
	mem[2487] = 4'b0000;
	mem[2488] = 4'b0000;
	mem[2489] = 4'b0000;
	mem[2490] = 4'b0000;
	mem[2491] = 4'b0000;
	mem[2492] = 4'b0000;
	mem[2493] = 4'b0000;
	mem[2494] = 4'b0000;
	mem[2495] = 4'b0000;
	mem[2496] = 4'b0000;
	mem[2497] = 4'b0000;
	mem[2498] = 4'b0000;
	mem[2499] = 4'b0000;
	mem[2500] = 4'b0001;
	mem[2501] = 4'b0000;
	mem[2502] = 4'b0000;
	mem[2503] = 4'b0000;
	mem[2504] = 4'b0000;
	mem[2505] = 4'b0000;
	mem[2506] = 4'b0000;
	mem[2507] = 4'b0000;
	mem[2508] = 4'b0000;
	mem[2509] = 4'b0000;
	mem[2510] = 4'b0000;
	mem[2511] = 4'b0000;
	mem[2512] = 4'b0000;
	mem[2513] = 4'b0000;
	mem[2514] = 4'b0000;
	mem[2515] = 4'b0000;
	mem[2516] = 4'b0000;
	mem[2517] = 4'b0000;
	mem[2518] = 4'b0000;
	mem[2519] = 4'b0000;
	mem[2520] = 4'b0000;
	mem[2521] = 4'b0000;
	mem[2522] = 4'b0000;
	mem[2523] = 4'b0000;
	mem[2524] = 4'b0000;
	mem[2525] = 4'b0000;
	mem[2526] = 4'b0000;
	mem[2527] = 4'b0000;
	mem[2528] = 4'b0000;
	mem[2529] = 4'b0000;
	mem[2530] = 4'b0000;
	mem[2531] = 4'b0000;
	mem[2532] = 4'b0000;
	mem[2533] = 4'b0000;
	mem[2534] = 4'b0000;
	mem[2535] = 4'b0000;
	mem[2536] = 4'b0000;
	mem[2537] = 4'b0000;
	mem[2538] = 4'b0000;
	mem[2539] = 4'b0000;
	mem[2540] = 4'b0000;
	mem[2541] = 4'b0000;
	mem[2542] = 4'b0000;
	mem[2543] = 4'b0000;
	mem[2544] = 4'b0000;
	mem[2545] = 4'b0000;
	mem[2546] = 4'b0000;
	mem[2547] = 4'b0000;
	mem[2548] = 4'b0000;
	mem[2549] = 4'b0000;
	mem[2550] = 4'b0000;
	mem[2551] = 4'b0000;
	mem[2552] = 4'b0000;
	mem[2553] = 4'b0000;
	mem[2554] = 4'b0000;
	mem[2555] = 4'b0000;
	mem[2556] = 4'b0000;
	mem[2557] = 4'b0000;
	mem[2558] = 4'b0000;
	mem[2559] = 4'b0000;
	mem[2560] = 4'b0000;
	mem[2561] = 4'b0000;
	mem[2562] = 4'b0000;
	mem[2563] = 4'b0000;
	mem[2564] = 4'b0000;
	mem[2565] = 4'b0000;
	mem[2566] = 4'b0000;
	mem[2567] = 4'b0000;
	mem[2568] = 4'b0000;
	mem[2569] = 4'b0000;
	mem[2570] = 4'b0000;
	mem[2571] = 4'b0000;
	mem[2572] = 4'b0000;
	mem[2573] = 4'b0000;
	mem[2574] = 4'b0000;
	mem[2575] = 4'b0000;
	mem[2576] = 4'b0000;
	mem[2577] = 4'b0000;
	mem[2578] = 4'b0000;
	mem[2579] = 4'b0001;
	mem[2580] = 4'b0001;
	mem[2581] = 4'b0001;
	mem[2582] = 4'b0001;
	mem[2583] = 4'b0001;
	mem[2584] = 4'b0001;
	mem[2585] = 4'b0000;
	mem[2586] = 4'b0000;
	mem[2587] = 4'b0000;
	mem[2588] = 4'b0000;
	mem[2589] = 4'b0000;
	mem[2590] = 4'b0000;
	mem[2591] = 4'b0000;
	mem[2592] = 4'b0000;
	mem[2593] = 4'b0000;
	mem[2594] = 4'b0000;
	mem[2595] = 4'b0000;
	mem[2596] = 4'b0000;
	mem[2597] = 4'b0000;
	mem[2598] = 4'b0000;
	mem[2599] = 4'b0000;
	mem[2600] = 4'b0000;
	mem[2601] = 4'b0000;
	mem[2602] = 4'b0000;
	mem[2603] = 4'b0000;
	mem[2604] = 4'b0000;
	mem[2605] = 4'b0000;
	mem[2606] = 4'b0000;
	mem[2607] = 4'b0000;
	mem[2608] = 4'b0000;
	mem[2609] = 4'b0000;
	mem[2610] = 4'b0000;
	mem[2611] = 4'b0000;
	mem[2612] = 4'b0000;
	mem[2613] = 4'b0000;
	mem[2614] = 4'b0000;
	mem[2615] = 4'b0000;
	mem[2616] = 4'b0000;
	mem[2617] = 4'b0000;
	mem[2618] = 4'b0000;
	mem[2619] = 4'b0000;
	mem[2620] = 4'b0000;
	mem[2621] = 4'b0000;
	mem[2622] = 4'b0000;
	mem[2623] = 4'b0000;
	mem[2624] = 4'b0000;
	mem[2625] = 4'b0000;
	mem[2626] = 4'b0000;
	mem[2627] = 4'b0001;
	mem[2628] = 4'b0001;
	mem[2629] = 4'b0000;
	mem[2630] = 4'b0000;
	mem[2631] = 4'b0000;
	mem[2632] = 4'b0000;
	mem[2633] = 4'b0000;
	mem[2634] = 4'b0000;
	mem[2635] = 4'b0000;
	mem[2636] = 4'b0000;
	mem[2637] = 4'b0000;
	mem[2638] = 4'b0000;
	mem[2639] = 4'b0000;
	mem[2640] = 4'b0000;
	mem[2641] = 4'b0000;
	mem[2642] = 4'b0000;
	mem[2643] = 4'b0000;
	mem[2644] = 4'b0000;
	mem[2645] = 4'b0000;
	mem[2646] = 4'b0000;
	mem[2647] = 4'b0000;
	mem[2648] = 4'b0000;
	mem[2649] = 4'b0000;
	mem[2650] = 4'b0000;
	mem[2651] = 4'b0000;
	mem[2652] = 4'b0000;
	mem[2653] = 4'b0000;
	mem[2654] = 4'b0000;
	mem[2655] = 4'b0000;
	mem[2656] = 4'b0000;
	mem[2657] = 4'b0000;
	mem[2658] = 4'b0000;
	mem[2659] = 4'b0000;
	mem[2660] = 4'b0000;
	mem[2661] = 4'b0000;
	mem[2662] = 4'b0000;
	mem[2663] = 4'b0000;
	mem[2664] = 4'b0000;
	mem[2665] = 4'b0000;
	mem[2666] = 4'b0000;
	mem[2667] = 4'b0000;
	mem[2668] = 4'b0000;
	mem[2669] = 4'b0000;
	mem[2670] = 4'b0000;
	mem[2671] = 4'b0000;
	mem[2672] = 4'b0000;
	mem[2673] = 4'b0000;
	mem[2674] = 4'b0000;
	mem[2675] = 4'b0000;
	mem[2676] = 4'b0000;
	mem[2677] = 4'b0000;
	mem[2678] = 4'b0000;
	mem[2679] = 4'b0000;
	mem[2680] = 4'b0000;
	mem[2681] = 4'b0000;
	mem[2682] = 4'b0000;
	mem[2683] = 4'b0000;
	mem[2684] = 4'b0000;
	mem[2685] = 4'b0000;
	mem[2686] = 4'b0000;
	mem[2687] = 4'b0000;
	mem[2688] = 4'b0000;
	mem[2689] = 4'b0000;
	mem[2690] = 4'b0000;
	mem[2691] = 4'b0000;
	mem[2692] = 4'b0000;
	mem[2693] = 4'b0000;
	mem[2694] = 4'b0000;
	mem[2695] = 4'b0000;
	mem[2696] = 4'b0000;
	mem[2697] = 4'b0000;
	mem[2698] = 4'b0000;
	mem[2699] = 4'b0000;
	mem[2700] = 4'b0000;
	mem[2701] = 4'b0000;
	mem[2702] = 4'b0000;
	mem[2703] = 4'b0000;
	mem[2704] = 4'b0000;
	mem[2705] = 4'b0000;
	mem[2706] = 4'b0000;
	mem[2707] = 4'b0000;
	mem[2708] = 4'b0000;
	mem[2709] = 4'b0000;
	mem[2710] = 4'b0000;
	mem[2711] = 4'b0000;
	mem[2712] = 4'b0000;
	mem[2713] = 4'b0000;
	mem[2714] = 4'b0000;
	mem[2715] = 4'b0000;
	mem[2716] = 4'b0000;
	mem[2717] = 4'b0000;
	mem[2718] = 4'b0000;
	mem[2719] = 4'b0000;
	mem[2720] = 4'b0000;
	mem[2721] = 4'b0000;
	mem[2722] = 4'b0000;
	mem[2723] = 4'b0000;
	mem[2724] = 4'b0000;
	mem[2725] = 4'b0000;
	mem[2726] = 4'b0000;
	mem[2727] = 4'b0000;
	mem[2728] = 4'b0000;
	mem[2729] = 4'b0000;
	mem[2730] = 4'b0000;
	mem[2731] = 4'b0000;
	mem[2732] = 4'b0000;
	mem[2733] = 4'b0000;
	mem[2734] = 4'b0000;
	mem[2735] = 4'b0000;
	mem[2736] = 4'b0000;
	mem[2737] = 4'b0000;
	mem[2738] = 4'b0000;
	mem[2739] = 4'b0000;
	mem[2740] = 4'b0000;
	mem[2741] = 4'b0000;
	mem[2742] = 4'b0000;
	mem[2743] = 4'b0000;
	mem[2744] = 4'b0000;
	mem[2745] = 4'b0000;
	mem[2746] = 4'b0000;
	mem[2747] = 4'b0000;
	mem[2748] = 4'b0000;
	mem[2749] = 4'b0000;
	mem[2750] = 4'b0001;
	mem[2751] = 4'b0000;
	mem[2752] = 4'b0000;
	mem[2753] = 4'b0000;
	mem[2754] = 4'b0001;
	mem[2755] = 4'b0001;
	mem[2756] = 4'b0000;
	mem[2757] = 4'b0000;
	mem[2758] = 4'b0000;
	mem[2759] = 4'b0000;
	mem[2760] = 4'b0000;
	mem[2761] = 4'b0000;
	mem[2762] = 4'b0000;
	mem[2763] = 4'b0000;
	mem[2764] = 4'b0000;
	mem[2765] = 4'b0000;
	mem[2766] = 4'b0000;
	mem[2767] = 4'b0000;
	mem[2768] = 4'b0000;
	mem[2769] = 4'b0000;
	mem[2770] = 4'b0000;
	mem[2771] = 4'b0000;
	mem[2772] = 4'b0000;
	mem[2773] = 4'b0000;
	mem[2774] = 4'b0000;
	mem[2775] = 4'b0000;
	mem[2776] = 4'b0000;
	mem[2777] = 4'b0000;
	mem[2778] = 4'b0000;
	mem[2779] = 4'b0000;
	mem[2780] = 4'b0000;
	mem[2781] = 4'b0000;
	mem[2782] = 4'b0000;
	mem[2783] = 4'b0000;
	mem[2784] = 4'b0000;
	mem[2785] = 4'b0000;
	mem[2786] = 4'b0000;
	mem[2787] = 4'b0000;
	mem[2788] = 4'b0000;
	mem[2789] = 4'b0000;
	mem[2790] = 4'b0000;
	mem[2791] = 4'b0000;
	mem[2792] = 4'b0000;
	mem[2793] = 4'b0000;
	mem[2794] = 4'b0000;
	mem[2795] = 4'b0000;
	mem[2796] = 4'b0000;
	mem[2797] = 4'b0000;
	mem[2798] = 4'b0000;
	mem[2799] = 4'b0000;
	mem[2800] = 4'b0000;
	mem[2801] = 4'b0000;
	mem[2802] = 4'b0000;
	mem[2803] = 4'b0000;
	mem[2804] = 4'b0000;
	mem[2805] = 4'b0000;
	mem[2806] = 4'b0000;
	mem[2807] = 4'b0000;
	mem[2808] = 4'b0000;
	mem[2809] = 4'b0000;
	mem[2810] = 4'b0000;
	mem[2811] = 4'b0000;
	mem[2812] = 4'b0000;
	mem[2813] = 4'b0000;
	mem[2814] = 4'b0000;
	mem[2815] = 4'b0000;
	mem[2816] = 4'b0000;
	mem[2817] = 4'b0000;
	mem[2818] = 4'b0000;
	mem[2819] = 4'b0000;
	mem[2820] = 4'b0000;
	mem[2821] = 4'b0000;
	mem[2822] = 4'b0000;
	mem[2823] = 4'b0000;
	mem[2824] = 4'b0000;
	mem[2825] = 4'b0000;
	mem[2826] = 4'b0000;
	mem[2827] = 4'b0000;
	mem[2828] = 4'b0000;
	mem[2829] = 4'b0000;
	mem[2830] = 4'b0000;
	mem[2831] = 4'b0000;
	mem[2832] = 4'b0000;
	mem[2833] = 4'b0000;
	mem[2834] = 4'b0000;
	mem[2835] = 4'b0000;
	mem[2836] = 4'b0000;
	mem[2837] = 4'b0000;
	mem[2838] = 4'b0000;
	mem[2839] = 4'b0000;
	mem[2840] = 4'b0000;
	mem[2841] = 4'b0000;
	mem[2842] = 4'b0000;
	mem[2843] = 4'b0000;
	mem[2844] = 4'b0000;
	mem[2845] = 4'b0000;
	mem[2846] = 4'b0000;
	mem[2847] = 4'b0000;
	mem[2848] = 4'b0000;
	mem[2849] = 4'b0000;
	mem[2850] = 4'b0000;
	mem[2851] = 4'b0000;
	mem[2852] = 4'b0000;
	mem[2853] = 4'b0000;
	mem[2854] = 4'b0000;
	mem[2855] = 4'b0000;
	mem[2856] = 4'b0000;
	mem[2857] = 4'b0000;
	mem[2858] = 4'b0000;
	mem[2859] = 4'b0000;
	mem[2860] = 4'b0000;
	mem[2861] = 4'b0000;
	mem[2862] = 4'b0000;
	mem[2863] = 4'b0000;
	mem[2864] = 4'b0000;
	mem[2865] = 4'b0000;
	mem[2866] = 4'b0000;
	mem[2867] = 4'b0000;
	mem[2868] = 4'b0000;
	mem[2869] = 4'b0000;
	mem[2870] = 4'b0000;
	mem[2871] = 4'b0000;
	mem[2872] = 4'b0000;
	mem[2873] = 4'b0000;
	mem[2874] = 4'b0000;
	mem[2875] = 4'b0000;
	mem[2876] = 4'b0000;
	mem[2877] = 4'b0000;
	mem[2878] = 4'b0000;
	mem[2879] = 4'b0000;
	mem[2880] = 4'b0001;
	mem[2881] = 4'b0001;
	mem[2882] = 4'b0000;
	mem[2883] = 4'b0000;
	mem[2884] = 4'b0000;
	mem[2885] = 4'b0000;
	mem[2886] = 4'b0000;
	mem[2887] = 4'b0000;
	mem[2888] = 4'b0000;
	mem[2889] = 4'b0000;
	mem[2890] = 4'b0000;
	mem[2891] = 4'b0000;
	mem[2892] = 4'b0000;
	mem[2893] = 4'b0000;
	mem[2894] = 4'b0000;
	mem[2895] = 4'b0000;
	mem[2896] = 4'b0000;
	mem[2897] = 4'b0000;
	mem[2898] = 4'b0000;
	mem[2899] = 4'b0000;
	mem[2900] = 4'b0000;
	mem[2901] = 4'b0000;
	mem[2902] = 4'b0000;
	mem[2903] = 4'b0000;
	mem[2904] = 4'b0000;
	mem[2905] = 4'b0000;
	mem[2906] = 4'b0000;
	mem[2907] = 4'b0000;
	mem[2908] = 4'b0000;
	mem[2909] = 4'b0000;
	mem[2910] = 4'b0000;
	mem[2911] = 4'b0000;
	mem[2912] = 4'b0000;
	mem[2913] = 4'b0000;
	mem[2914] = 4'b0000;
	mem[2915] = 4'b0000;
	mem[2916] = 4'b0000;
	mem[2917] = 4'b0000;
	mem[2918] = 4'b0000;
	mem[2919] = 4'b0000;
	mem[2920] = 4'b0000;
	mem[2921] = 4'b0000;
	mem[2922] = 4'b0000;
	mem[2923] = 4'b0000;
	mem[2924] = 4'b0000;
	mem[2925] = 4'b0000;
	mem[2926] = 4'b0000;
	mem[2927] = 4'b0000;
	mem[2928] = 4'b0000;
	mem[2929] = 4'b0000;
	mem[2930] = 4'b0000;
	mem[2931] = 4'b0000;
	mem[2932] = 4'b0000;
	mem[2933] = 4'b0000;
	mem[2934] = 4'b0000;
	mem[2935] = 4'b0000;
	mem[2936] = 4'b0000;
	mem[2937] = 4'b0000;
	mem[2938] = 4'b0000;
	mem[2939] = 4'b0000;
	mem[2940] = 4'b0000;
	mem[2941] = 4'b0000;
	mem[2942] = 4'b0000;
	mem[2943] = 4'b0000;
	mem[2944] = 4'b0000;
	mem[2945] = 4'b0000;
	mem[2946] = 4'b0000;
	mem[2947] = 4'b0000;
	mem[2948] = 4'b0000;
	mem[2949] = 4'b0000;
	mem[2950] = 4'b0000;
	mem[2951] = 4'b0000;
	mem[2952] = 4'b0000;
	mem[2953] = 4'b0000;
	mem[2954] = 4'b0000;
	mem[2955] = 4'b0000;
	mem[2956] = 4'b0000;
	mem[2957] = 4'b0000;
	mem[2958] = 4'b0000;
	mem[2959] = 4'b0000;
	mem[2960] = 4'b0000;
	mem[2961] = 4'b0000;
	mem[2962] = 4'b0000;
	mem[2963] = 4'b0000;
	mem[2964] = 4'b0000;
	mem[2965] = 4'b0000;
	mem[2966] = 4'b0000;
	mem[2967] = 4'b0000;
	mem[2968] = 4'b0000;
	mem[2969] = 4'b0000;
	mem[2970] = 4'b0000;
	mem[2971] = 4'b0000;
	mem[2972] = 4'b0000;
	mem[2973] = 4'b0000;
	mem[2974] = 4'b0000;
	mem[2975] = 4'b0000;
	mem[2976] = 4'b0000;
	mem[2977] = 4'b0000;
	mem[2978] = 4'b0000;
	mem[2979] = 4'b0000;
	mem[2980] = 4'b0000;
	mem[2981] = 4'b0000;
	mem[2982] = 4'b0000;
	mem[2983] = 4'b0000;
	mem[2984] = 4'b0000;
	mem[2985] = 4'b0000;
	mem[2986] = 4'b0000;
	mem[2987] = 4'b0000;
	mem[2988] = 4'b0000;
	mem[2989] = 4'b0000;
	mem[2990] = 4'b0000;
	mem[2991] = 4'b0000;
	mem[2992] = 4'b0000;
	mem[2993] = 4'b0000;
	mem[2994] = 4'b0000;
	mem[2995] = 4'b0000;
	mem[2996] = 4'b0000;
	mem[2997] = 4'b0000;
	mem[2998] = 4'b0000;
	mem[2999] = 4'b0000;
	mem[3000] = 4'b0000;
	mem[3001] = 4'b0000;
	mem[3002] = 4'b0000;
	mem[3003] = 4'b0000;
	mem[3004] = 4'b0000;
	mem[3005] = 4'b0000;
	mem[3006] = 4'b0000;
	mem[3007] = 4'b0000;
	mem[3008] = 4'b0000;
	mem[3009] = 4'b0000;
	mem[3010] = 4'b0000;
	mem[3011] = 4'b0000;
	mem[3012] = 4'b0000;
	mem[3013] = 4'b0000;
	mem[3014] = 4'b0000;
	mem[3015] = 4'b0000;
	mem[3016] = 4'b0000;
	mem[3017] = 4'b0000;
	mem[3018] = 4'b0000;
	mem[3019] = 4'b0000;
	mem[3020] = 4'b0000;
	mem[3021] = 4'b0000;
	mem[3022] = 4'b0000;
	mem[3023] = 4'b0000;
	mem[3024] = 4'b0000;
	mem[3025] = 4'b0000;
	mem[3026] = 4'b0000;
	mem[3027] = 4'b0000;
	mem[3028] = 4'b0000;
	mem[3029] = 4'b0000;
	mem[3030] = 4'b0000;
	mem[3031] = 4'b0000;
	mem[3032] = 4'b0000;
	mem[3033] = 4'b0000;
	mem[3034] = 4'b0000;
	mem[3035] = 4'b0000;
	mem[3036] = 4'b0000;
	mem[3037] = 4'b0000;
	mem[3038] = 4'b0000;
	mem[3039] = 4'b0000;
	mem[3040] = 4'b0000;
	mem[3041] = 4'b0000;
	mem[3042] = 4'b0000;
	mem[3043] = 4'b0000;
	mem[3044] = 4'b0000;
	mem[3045] = 4'b0000;
	mem[3046] = 4'b0000;
	mem[3047] = 4'b0000;
	mem[3048] = 4'b0000;
	mem[3049] = 4'b0000;
	mem[3050] = 4'b0000;
	mem[3051] = 4'b0000;
	mem[3052] = 4'b0000;
	mem[3053] = 4'b0000;
	mem[3054] = 4'b0000;
	mem[3055] = 4'b0000;
	mem[3056] = 4'b0000;
	mem[3057] = 4'b0000;
	mem[3058] = 4'b0000;
	mem[3059] = 4'b0000;
	mem[3060] = 4'b0000;
	mem[3061] = 4'b0000;
	mem[3062] = 4'b0000;
	mem[3063] = 4'b0000;
	mem[3064] = 4'b0000;
	mem[3065] = 4'b0000;
	mem[3066] = 4'b0000;
	mem[3067] = 4'b0000;
	mem[3068] = 4'b0000;
	mem[3069] = 4'b0000;
	mem[3070] = 4'b0000;
	mem[3071] = 4'b0000;
	mem[3072] = 4'b0000;
	mem[3073] = 4'b0000;
	mem[3074] = 4'b0000;
	mem[3075] = 4'b0000;
	mem[3076] = 4'b0000;
	mem[3077] = 4'b0000;
	mem[3078] = 4'b0000;
	mem[3079] = 4'b0000;
	mem[3080] = 4'b0000;
	mem[3081] = 4'b0000;
	mem[3082] = 4'b0000;
	mem[3083] = 4'b0000;
	mem[3084] = 4'b0000;
	mem[3085] = 4'b0000;
	mem[3086] = 4'b0000;
	mem[3087] = 4'b0000;
	mem[3088] = 4'b0000;
	mem[3089] = 4'b0000;
	mem[3090] = 4'b0000;
	mem[3091] = 4'b0000;
	mem[3092] = 4'b0000;
	mem[3093] = 4'b0000;
	mem[3094] = 4'b0000;
	mem[3095] = 4'b0000;
	mem[3096] = 4'b0000;
	mem[3097] = 4'b0000;
	mem[3098] = 4'b0000;
	mem[3099] = 4'b0000;
	mem[3100] = 4'b0000;
	mem[3101] = 4'b0000;
	mem[3102] = 4'b0000;
	mem[3103] = 4'b0000;
	mem[3104] = 4'b0000;
	mem[3105] = 4'b0000;
	mem[3106] = 4'b0000;
	mem[3107] = 4'b0000;
	mem[3108] = 4'b0000;
	mem[3109] = 4'b0000;
	mem[3110] = 4'b0000;
	mem[3111] = 4'b0000;
	mem[3112] = 4'b0000;
	mem[3113] = 4'b0000;
	mem[3114] = 4'b0000;
	mem[3115] = 4'b0000;
	mem[3116] = 4'b0000;
	mem[3117] = 4'b0000;
	mem[3118] = 4'b0000;
	mem[3119] = 4'b0000;
	mem[3120] = 4'b0000;
	mem[3121] = 4'b0000;
	mem[3122] = 4'b0000;
	mem[3123] = 4'b0000;
	mem[3124] = 4'b0000;
	mem[3125] = 4'b0000;
	mem[3126] = 4'b0000;
	mem[3127] = 4'b0000;
	mem[3128] = 4'b0000;
	mem[3129] = 4'b0000;
	mem[3130] = 4'b0000;
	mem[3131] = 4'b0000;
	mem[3132] = 4'b0000;
	mem[3133] = 4'b0000;
	mem[3134] = 4'b0000;
	mem[3135] = 4'b0000;
	mem[3136] = 4'b0000;
	mem[3137] = 4'b0000;
	mem[3138] = 4'b0000;
	mem[3139] = 4'b0000;
	mem[3140] = 4'b0000;
	mem[3141] = 4'b0000;
	mem[3142] = 4'b0000;
	mem[3143] = 4'b0000;
	mem[3144] = 4'b0000;
	mem[3145] = 4'b0000;
	mem[3146] = 4'b0000;
	mem[3147] = 4'b0000;
	mem[3148] = 4'b0000;
	mem[3149] = 4'b0000;
	mem[3150] = 4'b0000;
	mem[3151] = 4'b0000;
	mem[3152] = 4'b0000;
	mem[3153] = 4'b0000;
	mem[3154] = 4'b0000;
	mem[3155] = 4'b0000;
	mem[3156] = 4'b0000;
	mem[3157] = 4'b0000;
	mem[3158] = 4'b0000;
	mem[3159] = 4'b0000;
	mem[3160] = 4'b0000;
	mem[3161] = 4'b0000;
	mem[3162] = 4'b0000;
	mem[3163] = 4'b0000;
	mem[3164] = 4'b0000;
	mem[3165] = 4'b0000;
	mem[3166] = 4'b0000;
	mem[3167] = 4'b0000;
	mem[3168] = 4'b0000;
	mem[3169] = 4'b0000;
	mem[3170] = 4'b0000;
	mem[3171] = 4'b0000;
	mem[3172] = 4'b0000;
	mem[3173] = 4'b0000;
	mem[3174] = 4'b0000;
	mem[3175] = 4'b0000;
	mem[3176] = 4'b0000;
	mem[3177] = 4'b0000;
	mem[3178] = 4'b0000;
	mem[3179] = 4'b0000;
	mem[3180] = 4'b0000;
	mem[3181] = 4'b0000;
	mem[3182] = 4'b0000;
	mem[3183] = 4'b0000;
	mem[3184] = 4'b0000;
	mem[3185] = 4'b0000;
	mem[3186] = 4'b0000;
	mem[3187] = 4'b0000;
	mem[3188] = 4'b0000;
	mem[3189] = 4'b0000;
	mem[3190] = 4'b0000;
	mem[3191] = 4'b0000;
	mem[3192] = 4'b0000;
	mem[3193] = 4'b0000;
	mem[3194] = 4'b0000;
	mem[3195] = 4'b0000;
	mem[3196] = 4'b0000;
	mem[3197] = 4'b0000;
	mem[3198] = 4'b0000;
	mem[3199] = 4'b0000;
	mem[3200] = 4'b0000;
	mem[3201] = 4'b0000;
	mem[3202] = 4'b0000;
	mem[3203] = 4'b0000;
	mem[3204] = 4'b0000;
	mem[3205] = 4'b0000;
	mem[3206] = 4'b0000;
	mem[3207] = 4'b0000;
	mem[3208] = 4'b0000;
	mem[3209] = 4'b0000;
	mem[3210] = 4'b0000;
	mem[3211] = 4'b0000;
	mem[3212] = 4'b0000;
	mem[3213] = 4'b0000;
	mem[3214] = 4'b0000;
	mem[3215] = 4'b0000;
	mem[3216] = 4'b0000;
	mem[3217] = 4'b0000;
	mem[3218] = 4'b0000;
	mem[3219] = 4'b0000;
	mem[3220] = 4'b0000;
	mem[3221] = 4'b0000;
	mem[3222] = 4'b0000;
	mem[3223] = 4'b0000;
	mem[3224] = 4'b0000;
	mem[3225] = 4'b0000;
	mem[3226] = 4'b0000;
	mem[3227] = 4'b0000;
	mem[3228] = 4'b0000;
	mem[3229] = 4'b0000;
	mem[3230] = 4'b0000;
	mem[3231] = 4'b0000;
	mem[3232] = 4'b0000;
	mem[3233] = 4'b0000;
	mem[3234] = 4'b0000;
	mem[3235] = 4'b0000;
	mem[3236] = 4'b0000;
	mem[3237] = 4'b0000;
	mem[3238] = 4'b0000;
	mem[3239] = 4'b0000;
	mem[3240] = 4'b0000;
	mem[3241] = 4'b0000;
	mem[3242] = 4'b0000;
	mem[3243] = 4'b0000;
	mem[3244] = 4'b0000;
	mem[3245] = 4'b0000;
	mem[3246] = 4'b0000;
	mem[3247] = 4'b0000;
	mem[3248] = 4'b0000;
	mem[3249] = 4'b0000;
	mem[3250] = 4'b0000;
	mem[3251] = 4'b0000;
	mem[3252] = 4'b0000;
	mem[3253] = 4'b0000;
	mem[3254] = 4'b0000;
	mem[3255] = 4'b0000;
	mem[3256] = 4'b0000;
	mem[3257] = 4'b0000;
	mem[3258] = 4'b0000;
	mem[3259] = 4'b0000;
	mem[3260] = 4'b0000;
	mem[3261] = 4'b0000;
	mem[3262] = 4'b0001;
	mem[3263] = 4'b0000;
	mem[3264] = 4'b0000;
	mem[3265] = 4'b0000;
	mem[3266] = 4'b0000;
	mem[3267] = 4'b0000;
	mem[3268] = 4'b0000;
	mem[3269] = 4'b0000;
	mem[3270] = 4'b0000;
	mem[3271] = 4'b0000;
	mem[3272] = 4'b0000;
	mem[3273] = 4'b0000;
	mem[3274] = 4'b0000;
	mem[3275] = 4'b0000;
	mem[3276] = 4'b0000;
	mem[3277] = 4'b0000;
	mem[3278] = 4'b0000;
	mem[3279] = 4'b0000;
	mem[3280] = 4'b0000;
	mem[3281] = 4'b0000;
	mem[3282] = 4'b0000;
	mem[3283] = 4'b0000;
	mem[3284] = 4'b0000;
	mem[3285] = 4'b0000;
	mem[3286] = 4'b0000;
	mem[3287] = 4'b0000;
	mem[3288] = 4'b0000;
	mem[3289] = 4'b0000;
	mem[3290] = 4'b0000;
	mem[3291] = 4'b0000;
	mem[3292] = 4'b0000;
	mem[3293] = 4'b0000;
	mem[3294] = 4'b0000;
	mem[3295] = 4'b0000;
	mem[3296] = 4'b0000;
	mem[3297] = 4'b0000;
	mem[3298] = 4'b0000;
	mem[3299] = 4'b0000;
	mem[3300] = 4'b0000;
	mem[3301] = 4'b0000;
	mem[3302] = 4'b0000;
	mem[3303] = 4'b0000;
	mem[3304] = 4'b0000;
	mem[3305] = 4'b0000;
	mem[3306] = 4'b0000;
	mem[3307] = 4'b0000;
	mem[3308] = 4'b0000;
	mem[3309] = 4'b0000;
	mem[3310] = 4'b0000;
	mem[3311] = 4'b0000;
	mem[3312] = 4'b0000;
	mem[3313] = 4'b0000;
	mem[3314] = 4'b0000;
	mem[3315] = 4'b0000;
	mem[3316] = 4'b0000;
	mem[3317] = 4'b0000;
	mem[3318] = 4'b0000;
	mem[3319] = 4'b0000;
	mem[3320] = 4'b0000;
	mem[3321] = 4'b0000;
	mem[3322] = 4'b0000;
	mem[3323] = 4'b0000;
	mem[3324] = 4'b0000;
	mem[3325] = 4'b0000;
	mem[3326] = 4'b0000;
	mem[3327] = 4'b0000;
	mem[3328] = 4'b0000;
	mem[3329] = 4'b0000;
	mem[3330] = 4'b0000;
	mem[3331] = 4'b0000;
	mem[3332] = 4'b0000;
	mem[3333] = 4'b0000;
	mem[3334] = 4'b0000;
	mem[3335] = 4'b0000;
	mem[3336] = 4'b0000;
	mem[3337] = 4'b0000;
	mem[3338] = 4'b0000;
	mem[3339] = 4'b0000;
	mem[3340] = 4'b0000;
	mem[3341] = 4'b0000;
	mem[3342] = 4'b0000;
	mem[3343] = 4'b0000;
	mem[3344] = 4'b0000;
	mem[3345] = 4'b0000;
	mem[3346] = 4'b0001;
	mem[3347] = 4'b0001;
	mem[3348] = 4'b0000;
	mem[3349] = 4'b0000;
	mem[3350] = 4'b0000;
	mem[3351] = 4'b0000;
	mem[3352] = 4'b0000;
	mem[3353] = 4'b0000;
	mem[3354] = 4'b0000;
	mem[3355] = 4'b0000;
	mem[3356] = 4'b0000;
	mem[3357] = 4'b0000;
	mem[3358] = 4'b0000;
	mem[3359] = 4'b0000;
	mem[3360] = 4'b0000;
	mem[3361] = 4'b0000;
	mem[3362] = 4'b0000;
	mem[3363] = 4'b0000;
	mem[3364] = 4'b0000;
	mem[3365] = 4'b0000;
	mem[3366] = 4'b0000;
	mem[3367] = 4'b0000;
	mem[3368] = 4'b0000;
	mem[3369] = 4'b0000;
	mem[3370] = 4'b0000;
	mem[3371] = 4'b0000;
	mem[3372] = 4'b0000;
	mem[3373] = 4'b0000;
	mem[3374] = 4'b0000;
	mem[3375] = 4'b0000;
	mem[3376] = 4'b0000;
	mem[3377] = 4'b0000;
	mem[3378] = 4'b0000;
	mem[3379] = 4'b0000;
	mem[3380] = 4'b0000;
	mem[3381] = 4'b0000;
	mem[3382] = 4'b0000;
	mem[3383] = 4'b0000;
	mem[3384] = 4'b0000;
	mem[3385] = 4'b0000;
	mem[3386] = 4'b0000;
	mem[3387] = 4'b0000;
	mem[3388] = 4'b0000;
	mem[3389] = 4'b0001;
	mem[3390] = 4'b0001;
	mem[3391] = 4'b0000;
	mem[3392] = 4'b0000;
	mem[3393] = 4'b0000;
	mem[3394] = 4'b0000;
	mem[3395] = 4'b0000;
	mem[3396] = 4'b0000;
	mem[3397] = 4'b0000;
	mem[3398] = 4'b0000;
	mem[3399] = 4'b0000;
	mem[3400] = 4'b0000;
	mem[3401] = 4'b0000;
	mem[3402] = 4'b0000;
	mem[3403] = 4'b0000;
	mem[3404] = 4'b0000;
	mem[3405] = 4'b0000;
	mem[3406] = 4'b0000;
	mem[3407] = 4'b0000;
	mem[3408] = 4'b0000;
	mem[3409] = 4'b0000;
	mem[3410] = 4'b0000;
	mem[3411] = 4'b0000;
	mem[3412] = 4'b0000;
	mem[3413] = 4'b0000;
	mem[3414] = 4'b0000;
	mem[3415] = 4'b0000;
	mem[3416] = 4'b0000;
	mem[3417] = 4'b0000;
	mem[3418] = 4'b0000;
	mem[3419] = 4'b0000;
	mem[3420] = 4'b0000;
	mem[3421] = 4'b0000;
	mem[3422] = 4'b0000;
	mem[3423] = 4'b0000;
	mem[3424] = 4'b0000;
	mem[3425] = 4'b0000;
	mem[3426] = 4'b0000;
	mem[3427] = 4'b0000;
	mem[3428] = 4'b0000;
	mem[3429] = 4'b0000;
	mem[3430] = 4'b0000;
	mem[3431] = 4'b0000;
	mem[3432] = 4'b0000;
	mem[3433] = 4'b0000;
	mem[3434] = 4'b0000;
	mem[3435] = 4'b0000;
	mem[3436] = 4'b0000;
	mem[3437] = 4'b0000;
	mem[3438] = 4'b0000;
	mem[3439] = 4'b0000;
	mem[3440] = 4'b0000;
	mem[3441] = 4'b0000;
	mem[3442] = 4'b0000;
	mem[3443] = 4'b0000;
	mem[3444] = 4'b0000;
	mem[3445] = 4'b0000;
	mem[3446] = 4'b0000;
	mem[3447] = 4'b0000;
	mem[3448] = 4'b0000;
	mem[3449] = 4'b0000;
	mem[3450] = 4'b0000;
	mem[3451] = 4'b0000;
	mem[3452] = 4'b0000;
	mem[3453] = 4'b0000;
	mem[3454] = 4'b0000;
	mem[3455] = 4'b0000;
	mem[3456] = 4'b0000;
	mem[3457] = 4'b0000;
	mem[3458] = 4'b0000;
	mem[3459] = 4'b0000;
	mem[3460] = 4'b0000;
	mem[3461] = 4'b0000;
	mem[3462] = 4'b0000;
	mem[3463] = 4'b0000;
	mem[3464] = 4'b0000;
	mem[3465] = 4'b0000;
	mem[3466] = 4'b0000;
	mem[3467] = 4'b0000;
	mem[3468] = 4'b0000;
	mem[3469] = 4'b0000;
	mem[3470] = 4'b0000;
	mem[3471] = 4'b0000;
	mem[3472] = 4'b0000;
	mem[3473] = 4'b0001;
	mem[3474] = 4'b0001;
	mem[3475] = 4'b0000;
	mem[3476] = 4'b0000;
	mem[3477] = 4'b0000;
	mem[3478] = 4'b0000;
	mem[3479] = 4'b0000;
	mem[3480] = 4'b0000;
	mem[3481] = 4'b0000;
	mem[3482] = 4'b0000;
	mem[3483] = 4'b0000;
	mem[3484] = 4'b0000;
	mem[3485] = 4'b0000;
	mem[3486] = 4'b0000;
	mem[3487] = 4'b0000;
	mem[3488] = 4'b0000;
	mem[3489] = 4'b0000;
	mem[3490] = 4'b0000;
	mem[3491] = 4'b0000;
	mem[3492] = 4'b0000;
	mem[3493] = 4'b0000;
	mem[3494] = 4'b0000;
	mem[3495] = 4'b0000;
	mem[3496] = 4'b0000;
	mem[3497] = 4'b0000;
	mem[3498] = 4'b0000;
	mem[3499] = 4'b0000;
	mem[3500] = 4'b0000;
	mem[3501] = 4'b0000;
	mem[3502] = 4'b0000;
	mem[3503] = 4'b0000;
	mem[3504] = 4'b0000;
	mem[3505] = 4'b0000;
	mem[3506] = 4'b0000;
	mem[3507] = 4'b0000;
	mem[3508] = 4'b0000;
	mem[3509] = 4'b0000;
	mem[3510] = 4'b0000;
	mem[3511] = 4'b0000;
	mem[3512] = 4'b0000;
	mem[3513] = 4'b0000;
	mem[3514] = 4'b0000;
	mem[3515] = 4'b0000;
	mem[3516] = 4'b0000;
	mem[3517] = 4'b0000;
	mem[3518] = 4'b0000;
	mem[3519] = 4'b0000;
	mem[3520] = 4'b0000;
	mem[3521] = 4'b0000;
	mem[3522] = 4'b0000;
	mem[3523] = 4'b0000;
	mem[3524] = 4'b0000;
	mem[3525] = 4'b0000;
	mem[3526] = 4'b0000;
	mem[3527] = 4'b0000;
	mem[3528] = 4'b0000;
	mem[3529] = 4'b0000;
	mem[3530] = 4'b0000;
	mem[3531] = 4'b0000;
	mem[3532] = 4'b0000;
	mem[3533] = 4'b0000;
	mem[3534] = 4'b0000;
	mem[3535] = 4'b0000;
	mem[3536] = 4'b0000;
	mem[3537] = 4'b0000;
	mem[3538] = 4'b0000;
	mem[3539] = 4'b0000;
	mem[3540] = 4'b0000;
	mem[3541] = 4'b0000;
	mem[3542] = 4'b0000;
	mem[3543] = 4'b0000;
	mem[3544] = 4'b0000;
	mem[3545] = 4'b0000;
	mem[3546] = 4'b0000;
	mem[3547] = 4'b0000;
	mem[3548] = 4'b0000;
	mem[3549] = 4'b0000;
	mem[3550] = 4'b0000;
	mem[3551] = 4'b0000;
	mem[3552] = 4'b0000;
	mem[3553] = 4'b0000;
	mem[3554] = 4'b0000;
	mem[3555] = 4'b0000;
	mem[3556] = 4'b0000;
	mem[3557] = 4'b0000;
	mem[3558] = 4'b0000;
	mem[3559] = 4'b0000;
	mem[3560] = 4'b0000;
	mem[3561] = 4'b0000;
	mem[3562] = 4'b0000;
	mem[3563] = 4'b0000;
	mem[3564] = 4'b0000;
	mem[3565] = 4'b0000;
	mem[3566] = 4'b0000;
	mem[3567] = 4'b0000;
	mem[3568] = 4'b0000;
	mem[3569] = 4'b0000;
	mem[3570] = 4'b0000;
	mem[3571] = 4'b0000;
	mem[3572] = 4'b0000;
	mem[3573] = 4'b0000;
	mem[3574] = 4'b0000;
	mem[3575] = 4'b0000;
	mem[3576] = 4'b0000;
	mem[3577] = 4'b0000;
	mem[3578] = 4'b0000;
	mem[3579] = 4'b0000;
	mem[3580] = 4'b0000;
	mem[3581] = 4'b0000;
	mem[3582] = 4'b0000;
	mem[3583] = 4'b0000;
	mem[3584] = 4'b0000;
	mem[3585] = 4'b0000;
	mem[3586] = 4'b0000;
	mem[3587] = 4'b0000;
	mem[3588] = 4'b0000;
	mem[3589] = 4'b0000;
	mem[3590] = 4'b0000;
	mem[3591] = 4'b0000;
	mem[3592] = 4'b0000;
	mem[3593] = 4'b0000;
	mem[3594] = 4'b0000;
	mem[3595] = 4'b0000;
	mem[3596] = 4'b0000;
	mem[3597] = 4'b0000;
	mem[3598] = 4'b0000;
	mem[3599] = 4'b0000;
	mem[3600] = 4'b0001;
	mem[3601] = 4'b0001;
	mem[3602] = 4'b0000;
	mem[3603] = 4'b0000;
	mem[3604] = 4'b0000;
	mem[3605] = 4'b0000;
	mem[3606] = 4'b0000;
	mem[3607] = 4'b0000;
	mem[3608] = 4'b0000;
	mem[3609] = 4'b0000;
	mem[3610] = 4'b0000;
	mem[3611] = 4'b0000;
	mem[3612] = 4'b0000;
	mem[3613] = 4'b0000;
	mem[3614] = 4'b0000;
	mem[3615] = 4'b0000;
	mem[3616] = 4'b0000;
	mem[3617] = 4'b0000;
	mem[3618] = 4'b0000;
	mem[3619] = 4'b0000;
	mem[3620] = 4'b0000;
	mem[3621] = 4'b0000;
	mem[3622] = 4'b0000;
	mem[3623] = 4'b0000;
	mem[3624] = 4'b0000;
	mem[3625] = 4'b0000;
	mem[3626] = 4'b0000;
	mem[3627] = 4'b0000;
	mem[3628] = 4'b0000;
	mem[3629] = 4'b0000;
	mem[3630] = 4'b0000;
	mem[3631] = 4'b0000;
	mem[3632] = 4'b0000;
	mem[3633] = 4'b0000;
	mem[3634] = 4'b0000;
	mem[3635] = 4'b0000;
	mem[3636] = 4'b0000;
	mem[3637] = 4'b0000;
	mem[3638] = 4'b0000;
	mem[3639] = 4'b0000;
	mem[3640] = 4'b0000;
	mem[3641] = 4'b0000;
	mem[3642] = 4'b0000;
	mem[3643] = 4'b0000;
	mem[3644] = 4'b0000;
	mem[3645] = 4'b0000;
	mem[3646] = 4'b0000;
	mem[3647] = 4'b0000;
	mem[3648] = 4'b0000;
	mem[3649] = 4'b0000;
	mem[3650] = 4'b0000;
	mem[3651] = 4'b0000;
	mem[3652] = 4'b0000;
	mem[3653] = 4'b0000;
	mem[3654] = 4'b0000;
	mem[3655] = 4'b0000;
	mem[3656] = 4'b0000;
	mem[3657] = 4'b0000;
	mem[3658] = 4'b0000;
	mem[3659] = 4'b0000;
	mem[3660] = 4'b0000;
	mem[3661] = 4'b0000;
	mem[3662] = 4'b0000;
	mem[3663] = 4'b0000;
	mem[3664] = 4'b0000;
	mem[3665] = 4'b0000;
	mem[3666] = 4'b0000;
	mem[3667] = 4'b0000;
	mem[3668] = 4'b0000;
	mem[3669] = 4'b0000;
	mem[3670] = 4'b0000;
	mem[3671] = 4'b0000;
	mem[3672] = 4'b0000;
	mem[3673] = 4'b0000;
	mem[3674] = 4'b0000;
	mem[3675] = 4'b0000;
	mem[3676] = 4'b0000;
	mem[3677] = 4'b0000;
	mem[3678] = 4'b0000;
	mem[3679] = 4'b0000;
	mem[3680] = 4'b0000;
	mem[3681] = 4'b0000;
	mem[3682] = 4'b0000;
	mem[3683] = 4'b0000;
	mem[3684] = 4'b0000;
	mem[3685] = 4'b0000;
	mem[3686] = 4'b0000;
	mem[3687] = 4'b0000;
	mem[3688] = 4'b0000;
	mem[3689] = 4'b0000;
	mem[3690] = 4'b0000;
	mem[3691] = 4'b0000;
	mem[3692] = 4'b0000;
	mem[3693] = 4'b0000;
	mem[3694] = 4'b0000;
	mem[3695] = 4'b0000;
	mem[3696] = 4'b0000;
	mem[3697] = 4'b0000;
	mem[3698] = 4'b0000;
	mem[3699] = 4'b0000;
	mem[3700] = 4'b0000;
	mem[3701] = 4'b0000;
	mem[3702] = 4'b0000;
	mem[3703] = 4'b0000;
	mem[3704] = 4'b0000;
	mem[3705] = 4'b0000;
	mem[3706] = 4'b0000;
	mem[3707] = 4'b0000;
	mem[3708] = 4'b0000;
	mem[3709] = 4'b0000;
	mem[3710] = 4'b0000;
	mem[3711] = 4'b0000;
	mem[3712] = 4'b0000;
	mem[3713] = 4'b0000;
	mem[3714] = 4'b0000;
	mem[3715] = 4'b0000;
	mem[3716] = 4'b0000;
	mem[3717] = 4'b0000;
	mem[3718] = 4'b0000;
	mem[3719] = 4'b0000;
	mem[3720] = 4'b0000;
	mem[3721] = 4'b0000;
	mem[3722] = 4'b0000;
	mem[3723] = 4'b0000;
	mem[3724] = 4'b0000;
	mem[3725] = 4'b0000;
	mem[3726] = 4'b0000;
	mem[3727] = 4'b0000;
	mem[3728] = 4'b0000;
	mem[3729] = 4'b0000;
	mem[3730] = 4'b0000;
	mem[3731] = 4'b0000;
	mem[3732] = 4'b0000;
	mem[3733] = 4'b0000;
	mem[3734] = 4'b0000;
	mem[3735] = 4'b0000;
	mem[3736] = 4'b0000;
	mem[3737] = 4'b0000;
	mem[3738] = 4'b0000;
	mem[3739] = 4'b0000;
	mem[3740] = 4'b0000;
	mem[3741] = 4'b0000;
	mem[3742] = 4'b0000;
	mem[3743] = 4'b0000;
	mem[3744] = 4'b0000;
	mem[3745] = 4'b0000;
	mem[3746] = 4'b0000;
	mem[3747] = 4'b0000;
	mem[3748] = 4'b0000;
	mem[3749] = 4'b0000;
	mem[3750] = 4'b0000;
	mem[3751] = 4'b0000;
	mem[3752] = 4'b0000;
	mem[3753] = 4'b0000;
	mem[3754] = 4'b0000;
	mem[3755] = 4'b0000;
	mem[3756] = 4'b0000;
	mem[3757] = 4'b0000;
	mem[3758] = 4'b0000;
	mem[3759] = 4'b0000;
	mem[3760] = 4'b0000;
	mem[3761] = 4'b0000;
	mem[3762] = 4'b0000;
	mem[3763] = 4'b0000;
	mem[3764] = 4'b0000;
	mem[3765] = 4'b0000;
	mem[3766] = 4'b0000;
	mem[3767] = 4'b0000;
	mem[3768] = 4'b0000;
	mem[3769] = 4'b0000;
	mem[3770] = 4'b0000;
	mem[3771] = 4'b0000;
	mem[3772] = 4'b0000;
	mem[3773] = 4'b0000;
	mem[3774] = 4'b0000;
	mem[3775] = 4'b0000;
	mem[3776] = 4'b0000;
	mem[3777] = 4'b0000;
	mem[3778] = 4'b0000;
	mem[3779] = 4'b0000;
	mem[3780] = 4'b0000;
	mem[3781] = 4'b0000;
	mem[3782] = 4'b0000;
	mem[3783] = 4'b0000;
	mem[3784] = 4'b0000;
	mem[3785] = 4'b0000;
	mem[3786] = 4'b0000;
	mem[3787] = 4'b0000;
	mem[3788] = 4'b0000;
	mem[3789] = 4'b0000;
	mem[3790] = 4'b0000;
	mem[3791] = 4'b0000;
	mem[3792] = 4'b0000;
	mem[3793] = 4'b0000;
	mem[3794] = 4'b0000;
	mem[3795] = 4'b0000;
	mem[3796] = 4'b0000;
	mem[3797] = 4'b0000;
	mem[3798] = 4'b0000;
	mem[3799] = 4'b0000;
	mem[3800] = 4'b0000;
	mem[3801] = 4'b0000;
	mem[3802] = 4'b0000;
	mem[3803] = 4'b0000;
	mem[3804] = 4'b0000;
	mem[3805] = 4'b0000;
	mem[3806] = 4'b0000;
	mem[3807] = 4'b0000;
	mem[3808] = 4'b0000;
	mem[3809] = 4'b0000;
	mem[3810] = 4'b0000;
	mem[3811] = 4'b0000;
	mem[3812] = 4'b0000;
	mem[3813] = 4'b0000;
	mem[3814] = 4'b0000;
	mem[3815] = 4'b0000;
	mem[3816] = 4'b0000;
	mem[3817] = 4'b0000;
	mem[3818] = 4'b0000;
	mem[3819] = 4'b0000;
	mem[3820] = 4'b0000;
	mem[3821] = 4'b0000;
	mem[3822] = 4'b0000;
	mem[3823] = 4'b0000;
	mem[3824] = 4'b0000;
	mem[3825] = 4'b0000;
	mem[3826] = 4'b0000;
	mem[3827] = 4'b0000;
	mem[3828] = 4'b0000;
	mem[3829] = 4'b0000;
	mem[3830] = 4'b0000;
	mem[3831] = 4'b0000;
	mem[3832] = 4'b0000;
	mem[3833] = 4'b0000;
	mem[3834] = 4'b0000;
	mem[3835] = 4'b0000;
	mem[3836] = 4'b0000;
	mem[3837] = 4'b0000;
	mem[3838] = 4'b0000;
	mem[3839] = 4'b0000;
	mem[3840] = 4'b0000;
	mem[3841] = 4'b0000;
	mem[3842] = 4'b0000;
	mem[3843] = 4'b0000;
	mem[3844] = 4'b0000;
	mem[3845] = 4'b0000;
	mem[3846] = 4'b0000;
	mem[3847] = 4'b0000;
	mem[3848] = 4'b0000;
	mem[3849] = 4'b0000;
	mem[3850] = 4'b0000;
	mem[3851] = 4'b0000;
	mem[3852] = 4'b0000;
	mem[3853] = 4'b0000;
	mem[3854] = 4'b0000;
	mem[3855] = 4'b0000;
	mem[3856] = 4'b0000;
	mem[3857] = 4'b0000;
	mem[3858] = 4'b0000;
	mem[3859] = 4'b0000;
	mem[3860] = 4'b0000;
	mem[3861] = 4'b0000;
	mem[3862] = 4'b0000;
	mem[3863] = 4'b0000;
	mem[3864] = 4'b0000;
	mem[3865] = 4'b0000;
	mem[3866] = 4'b0000;
	mem[3867] = 4'b0000;
	mem[3868] = 4'b0000;
	mem[3869] = 4'b0000;
	mem[3870] = 4'b0000;
	mem[3871] = 4'b0000;
	mem[3872] = 4'b0000;
	mem[3873] = 4'b0000;
	mem[3874] = 4'b0000;
	mem[3875] = 4'b0000;
	mem[3876] = 4'b0000;
	mem[3877] = 4'b0000;
	mem[3878] = 4'b0000;
	mem[3879] = 4'b0000;
	mem[3880] = 4'b0000;
	mem[3881] = 4'b0000;
	mem[3882] = 4'b0000;
	mem[3883] = 4'b0000;
	mem[3884] = 4'b0000;
	mem[3885] = 4'b0000;
	mem[3886] = 4'b0000;
	mem[3887] = 4'b0000;
	mem[3888] = 4'b0000;
	mem[3889] = 4'b0000;
	mem[3890] = 4'b0000;
	mem[3891] = 4'b0000;
	mem[3892] = 4'b0000;
	mem[3893] = 4'b0000;
	mem[3894] = 4'b0000;
	mem[3895] = 4'b0000;
	mem[3896] = 4'b0000;
	mem[3897] = 4'b0000;
	mem[3898] = 4'b0000;
	mem[3899] = 4'b0000;
	mem[3900] = 4'b0000;
	mem[3901] = 4'b0000;
	mem[3902] = 4'b0000;
	mem[3903] = 4'b0000;
	mem[3904] = 4'b0000;
	mem[3905] = 4'b0000;
	mem[3906] = 4'b0000;
	mem[3907] = 4'b0000;
	mem[3908] = 4'b0000;
	mem[3909] = 4'b0000;
	mem[3910] = 4'b0000;
	mem[3911] = 4'b0000;
	mem[3912] = 4'b0000;
	mem[3913] = 4'b0000;
	mem[3914] = 4'b0000;
	mem[3915] = 4'b0000;
	mem[3916] = 4'b0000;
	mem[3917] = 4'b0000;
	mem[3918] = 4'b0000;
	mem[3919] = 4'b0000;
	mem[3920] = 4'b0000;
	mem[3921] = 4'b0000;
	mem[3922] = 4'b0000;
	mem[3923] = 4'b0000;
	mem[3924] = 4'b0000;
	mem[3925] = 4'b0000;
	mem[3926] = 4'b0000;
	mem[3927] = 4'b0000;
	mem[3928] = 4'b0000;
	mem[3929] = 4'b0000;
	mem[3930] = 4'b0000;
	mem[3931] = 4'b0000;
	mem[3932] = 4'b0000;
	mem[3933] = 4'b0000;
	mem[3934] = 4'b0000;
	mem[3935] = 4'b0000;
	mem[3936] = 4'b0000;
	mem[3937] = 4'b0000;
	mem[3938] = 4'b0000;
	mem[3939] = 4'b0000;
	mem[3940] = 4'b0000;
	mem[3941] = 4'b0000;
	mem[3942] = 4'b0000;
	mem[3943] = 4'b0000;
	mem[3944] = 4'b0000;
	mem[3945] = 4'b0000;
	mem[3946] = 4'b0000;
	mem[3947] = 4'b0000;
	mem[3948] = 4'b0000;
	mem[3949] = 4'b0000;
	mem[3950] = 4'b0000;
	mem[3951] = 4'b0000;
	mem[3952] = 4'b0000;
	mem[3953] = 4'b0000;
	mem[3954] = 4'b0000;
	mem[3955] = 4'b0000;
	mem[3956] = 4'b0000;
	mem[3957] = 4'b0000;
	mem[3958] = 4'b0000;
	mem[3959] = 4'b0000;
	mem[3960] = 4'b0000;
	mem[3961] = 4'b0000;
	mem[3962] = 4'b0000;
	mem[3963] = 4'b0000;
	mem[3964] = 4'b0000;
	mem[3965] = 4'b0000;
	mem[3966] = 4'b0000;
	mem[3967] = 4'b0000;
	mem[3968] = 4'b0000;
	mem[3969] = 4'b0000;
	mem[3970] = 4'b0000;
	mem[3971] = 4'b0000;
	mem[3972] = 4'b0000;
	mem[3973] = 4'b0000;
	mem[3974] = 4'b0000;
	mem[3975] = 4'b0000;
	mem[3976] = 4'b0000;
	mem[3977] = 4'b0000;
	mem[3978] = 4'b0000;
	mem[3979] = 4'b0000;
	mem[3980] = 4'b0000;
	mem[3981] = 4'b0000;
	mem[3982] = 4'b0000;
	mem[3983] = 4'b0000;
	mem[3984] = 4'b0000;
	mem[3985] = 4'b0000;
	mem[3986] = 4'b0000;
	mem[3987] = 4'b0000;
	mem[3988] = 4'b0000;
	mem[3989] = 4'b0000;
	mem[3990] = 4'b0000;
	mem[3991] = 4'b0000;
	mem[3992] = 4'b0000;
	mem[3993] = 4'b0000;
	mem[3994] = 4'b0000;
	mem[3995] = 4'b0000;
	mem[3996] = 4'b0000;
	mem[3997] = 4'b0000;
	mem[3998] = 4'b0000;
	mem[3999] = 4'b0000;
	mem[4000] = 4'b0000;
	mem[4001] = 4'b0000;
	mem[4002] = 4'b0000;
	mem[4003] = 4'b0000;
	mem[4004] = 4'b0000;
	mem[4005] = 4'b0000;
	mem[4006] = 4'b0000;
	mem[4007] = 4'b0000;
	mem[4008] = 4'b0000;
	mem[4009] = 4'b0000;
	mem[4010] = 4'b0000;
	mem[4011] = 4'b0000;
	mem[4012] = 4'b0000;
	mem[4013] = 4'b0000;
	mem[4014] = 4'b0000;
	mem[4015] = 4'b0000;
	mem[4016] = 4'b0000;
	mem[4017] = 4'b0000;
	mem[4018] = 4'b0000;
	mem[4019] = 4'b0000;
	mem[4020] = 4'b0000;
	mem[4021] = 4'b0000;
	mem[4022] = 4'b0000;
	mem[4023] = 4'b0000;
	mem[4024] = 4'b0000;
	mem[4025] = 4'b0000;
	mem[4026] = 4'b0000;
	mem[4027] = 4'b0000;
	mem[4028] = 4'b0000;
	mem[4029] = 4'b0000;
	mem[4030] = 4'b0000;
	mem[4031] = 4'b0000;
	mem[4032] = 4'b0000;
	mem[4033] = 4'b0000;
	mem[4034] = 4'b0000;
	mem[4035] = 4'b0000;
	mem[4036] = 4'b0000;
	mem[4037] = 4'b0000;
	mem[4038] = 4'b0000;
	mem[4039] = 4'b0000;
	mem[4040] = 4'b0000;
	mem[4041] = 4'b0000;
	mem[4042] = 4'b0000;
	mem[4043] = 4'b0000;
	mem[4044] = 4'b0000;
	mem[4045] = 4'b0000;
	mem[4046] = 4'b0000;
	mem[4047] = 4'b0000;
	mem[4048] = 4'b0000;
	mem[4049] = 4'b0000;
	mem[4050] = 4'b0000;
	mem[4051] = 4'b0000;
	mem[4052] = 4'b0000;
	mem[4053] = 4'b0000;
	mem[4054] = 4'b0000;
	mem[4055] = 4'b0000;
	mem[4056] = 4'b0000;
	mem[4057] = 4'b0000;
	mem[4058] = 4'b0000;
	mem[4059] = 4'b0000;
	mem[4060] = 4'b0000;
	mem[4061] = 4'b0000;
	mem[4062] = 4'b0000;
	mem[4063] = 4'b0000;
	mem[4064] = 4'b0000;
	mem[4065] = 4'b0000;
	mem[4066] = 4'b0000;
	mem[4067] = 4'b0000;
	mem[4068] = 4'b0000;
	mem[4069] = 4'b0000;
	mem[4070] = 4'b0000;
	mem[4071] = 4'b0000;
	mem[4072] = 4'b0000;
	mem[4073] = 4'b0000;
	mem[4074] = 4'b0000;
	mem[4075] = 4'b0000;
	mem[4076] = 4'b0000;
	mem[4077] = 4'b0000;
	mem[4078] = 4'b0000;
	mem[4079] = 4'b0000;
	mem[4080] = 4'b0000;
	mem[4081] = 4'b0000;
	mem[4082] = 4'b0000;
	mem[4083] = 4'b0000;
	mem[4084] = 4'b0000;
	mem[4085] = 4'b0000;
	mem[4086] = 4'b0000;
	mem[4087] = 4'b0000;
	mem[4088] = 4'b0000;
	mem[4089] = 4'b0000;
	mem[4090] = 4'b0000;
	mem[4091] = 4'b0000;
	mem[4092] = 4'b0000;
	mem[4093] = 4'b0000;
	mem[4094] = 4'b0000;
	mem[4095] = 4'b0000;
end
endmodule

